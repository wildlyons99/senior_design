library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;entity background_rom is    port(
        clk : in std_logic;
        xadr: in unsigned(1 downto 0);
        yadr : in unsigned(1 downto 0); -- 0-1023
        grayScale : out std_logic_vector(7 downto 0)
        );
end background_rom;

architecture synth of background_rom is
signal totaladr : std_logic_vector(3 downto 0);
begin
    process (clk) begin
        if rising_edge(clk) then
            case totaladr is
                when "0000" => rgb <= "00000000";
                when "0001" => rgb <= "00000000";
                when "0010" => rgb <= "00000000";
                when "0011" => rgb <= "00000000";
                when "0100" => rgb <= "00000000";
                when "0101" => rgb <= "00000000";
                when "0110" => rgb <= "00000000";
                when "0111" => rgb <= "00000000";
                when "1000" => rgb <= "00000000";
                when "1001" => rgb <= "00000000";
                when "1010" => rgb <= "00000000";
                when "1011" => rgb <= "00000000";
                when "1100" => rgb <= "00000000";
                when "1101" => rgb <= "00000000";
                when "1110" => rgb <= "00000000";
                when "1111" => rgb <= "00000000";
                when "10000" => rgb <= "00000000";
                when "10001" => rgb <= "00000000";
                when "10010" => rgb <= "00000000";
                when "10011" => rgb <= "00000000";
                when "10100" => rgb <= "00000000";
                when "10101" => rgb <= "00000000";
                when "10110" => rgb <= "00000000";
                when "10111" => rgb <= "00000000";
                when "11000" => rgb <= "00000000";
                when "11001" => rgb <= "00000000";
                when "11010" => rgb <= "00000000";
                when "11011" => rgb <= "00000000";
                when "11100" => rgb <= "00000000";
                when "11101" => rgb <= "00000000";
                when "11110" => rgb <= "00000000";
                when "11111" => rgb <= "00000000";
                when "100000" => rgb <= "00000000";
                when "100001" => rgb <= "00000000";
                when "100010" => rgb <= "00000000";
                when "100011" => rgb <= "00000000";
                when "100100" => rgb <= "00000000";
                when "100101" => rgb <= "00000000";
                when "100110" => rgb <= "00000000";
                when "100111" => rgb <= "00000000";
                when "101000" => rgb <= "00000000";
                when "101001" => rgb <= "00000000";
                when "101010" => rgb <= "00000000";
                when "101011" => rgb <= "00000000";
                when "101100" => rgb <= "00000000";
                when "101101" => rgb <= "00000000";
                when "101110" => rgb <= "00000000";
                when "101111" => rgb <= "00000000";
                when "110000" => rgb <= "00000000";
                when "110001" => rgb <= "00000000";
                when "110010" => rgb <= "00000000";
                when "110011" => rgb <= "00000000";
                when "110100" => rgb <= "00000000";
                when "110101" => rgb <= "00000000";
                when "110110" => rgb <= "00000000";
                when "110111" => rgb <= "00000000";
                when "111000" => rgb <= "00000000";
                when "111001" => rgb <= "00000000";
                when "111010" => rgb <= "00000000";
                when "111011" => rgb <= "00000000";
                when "111100" => rgb <= "00000000";
                when "111101" => rgb <= "00000000";
                when "111110" => rgb <= "00000000";
                when "111111" => rgb <= "00000000";
                when "1000000" => rgb <= "00000000";
                when "1000001" => rgb <= "00000000";
                when "1000010" => rgb <= "00000000";
                when "1000011" => rgb <= "00000000";
                when "1000100" => rgb <= "00000000";
                when "1000101" => rgb <= "00000000";
                when "1000110" => rgb <= "00000000";
                when "1000111" => rgb <= "00000000";
                when "1001000" => rgb <= "00000000";
                when "1001001" => rgb <= "00000000";
                when "1001010" => rgb <= "00000000";
                when "1001011" => rgb <= "00000000";
                when "1001100" => rgb <= "00000000";
                when "1001101" => rgb <= "00000000";
                when "1001110" => rgb <= "00000000";
                when "1001111" => rgb <= "00000000";
                when "1010000" => rgb <= "00000000";
                when "1010001" => rgb <= "00000000";
                when "1010010" => rgb <= "00000000";
                when "1010011" => rgb <= "00000000";
                when "1010100" => rgb <= "00000000";
                when "1010101" => rgb <= "00000000";
                when "1010110" => rgb <= "00000000";
                when "1010111" => rgb <= "00000000";
                when "1011000" => rgb <= "00000000";
                when "1011001" => rgb <= "00000000";
                when "1011010" => rgb <= "00000000";
                when "1011011" => rgb <= "00000000";
                when "1011100" => rgb <= "00000000";
                when "1011101" => rgb <= "00000000";
                when "1011110" => rgb <= "00000000";
                when "1011111" => rgb <= "00000000";
                when "1100000" => rgb <= "00000000";
                when "1100001" => rgb <= "00000000";
                when "1100010" => rgb <= "00000000";
                when "1100011" => rgb <= "00000000";
                when "1100100" => rgb <= "00000000";
                when "1100101" => rgb <= "00000000";
                when "1100110" => rgb <= "00000000";
                when "1100111" => rgb <= "00000000";
                when "1101000" => rgb <= "00000000";
                when "1101001" => rgb <= "00000000";
                when "1101010" => rgb <= "00000000";
                when "1101011" => rgb <= "00000000";
                when "1101100" => rgb <= "00000000";
                when "1101101" => rgb <= "00000000";
                when "1101110" => rgb <= "00000000";
                when "1101111" => rgb <= "00000000";
                when "1110000" => rgb <= "00000000";
                when "1110001" => rgb <= "00000000";
                when "1110010" => rgb <= "00000000";
                when "1110011" => rgb <= "00000000";
                when "1110100" => rgb <= "00000000";
                when "1110101" => rgb <= "00000000";
                when "1110110" => rgb <= "00000000";
                when "1110111" => rgb <= "00000000";
                when "1111000" => rgb <= "00000000";
                when "1111001" => rgb <= "00000000";
                when "1111010" => rgb <= "00000000";
                when "1111011" => rgb <= "01101001";
                when "1111100" => rgb <= "11100011";
                when "1111101" => rgb <= "01111100";
                when "1111110" => rgb <= "10110110";
                when "1111111" => rgb <= "01111001";
                when "10000000" => rgb <= "00000000";
                when "10000001" => rgb <= "00000000";
                when "10000010" => rgb <= "00000000";
                when "10000011" => rgb <= "00000000";
                when "10000100" => rgb <= "00000000";
                when "10000101" => rgb <= "00000000";
                when "10000110" => rgb <= "00000000";
                when "10000111" => rgb <= "00000000";
                when "10001000" => rgb <= "00000000";
                when "10001001" => rgb <= "00000000";
                when "10001010" => rgb <= "00000000";
                when "10001011" => rgb <= "00000000";
                when "10001100" => rgb <= "00000000";
                when "10001101" => rgb <= "00000000";
                when "10001110" => rgb <= "00000000";
                when "10001111" => rgb <= "00000000";
                when "10010000" => rgb <= "00000000";
                when "10010001" => rgb <= "00000000";
                when "10010010" => rgb <= "00000000";
                when "10010011" => rgb <= "00000000";
                when "10010100" => rgb <= "00000000";
                when "10010101" => rgb <= "00000000";
                when "10010110" => rgb <= "00010011";
                when "10010111" => rgb <= "11111000";
                when "10011000" => rgb <= "11111110";
                when "10011001" => rgb <= "11111101";
                when "10011010" => rgb <= "11111110";
                when "10011011" => rgb <= "11111110";
                when "10011100" => rgb <= "01111101";
                when "10011101" => rgb <= "00000000";
                when "10011110" => rgb <= "00000000";
                when "10011111" => rgb <= "00000000";
                when "10100000" => rgb <= "00000000";
                when "10100001" => rgb <= "00000000";
                when "10100010" => rgb <= "00000000";
                when "10100011" => rgb <= "00000000";
                when "10100100" => rgb <= "00000000";
                when "10100101" => rgb <= "00000000";
                when "10100110" => rgb <= "00000000";
                when "10100111" => rgb <= "00000000";
                when "10101000" => rgb <= "00000000";
                when "10101001" => rgb <= "00000000";
                when "10101010" => rgb <= "00000000";
                when "10101011" => rgb <= "00000000";
                when "10101100" => rgb <= "00000000";
                when "10101101" => rgb <= "00000000";
                when "10101110" => rgb <= "00000000";
                when "10101111" => rgb <= "00000000";
                when "10110000" => rgb <= "00000000";
                when "10110001" => rgb <= "00000000";
                when "10110010" => rgb <= "01001100";
                when "10110011" => rgb <= "11111110";
                when "10110100" => rgb <= "10101100";
                when "10110101" => rgb <= "01011110";
                when "10110110" => rgb <= "10100110";
                when "10110111" => rgb <= "11111000";
                when "10111000" => rgb <= "11110100";
                when "10111001" => rgb <= "01000100";
                when "10111010" => rgb <= "00000000";
                when "10111011" => rgb <= "00000000";
                when "10111100" => rgb <= "00000000";
                when "10111101" => rgb <= "00000000";
                when "10111110" => rgb <= "00000000";
                when "10111111" => rgb <= "00000000";
                when "11000000" => rgb <= "00000000";
                when "11000001" => rgb <= "00000000";
                when "11000010" => rgb <= "00000000";
                when "11000011" => rgb <= "00000000";
                when "11000100" => rgb <= "00000000";
                when "11000101" => rgb <= "00000000";
                when "11000110" => rgb <= "00000000";
                when "11000111" => rgb <= "00000000";
                when "11001000" => rgb <= "00000000";
                when "11001001" => rgb <= "00000000";
                when "11001010" => rgb <= "00000000";
                when "11001011" => rgb <= "00000000";
                when "11001100" => rgb <= "00000000";
                when "11001101" => rgb <= "00000000";
                when "11001110" => rgb <= "11001011";
                when "11001111" => rgb <= "11111110";
                when "11010000" => rgb <= "01000001";
                when "11010001" => rgb <= "00000000";
                when "11010010" => rgb <= "00000000";
                when "11010011" => rgb <= "01010110";
                when "11010100" => rgb <= "11111110";
                when "11010101" => rgb <= "11011100";
                when "11010110" => rgb <= "00011001";
                when "11010111" => rgb <= "00000000";
                when "11011000" => rgb <= "00000000";
                when "11011001" => rgb <= "00000000";
                when "11011010" => rgb <= "00000000";
                when "11011011" => rgb <= "00000000";
                when "11011100" => rgb <= "00000000";
                when "11011101" => rgb <= "00000000";
                when "11011110" => rgb <= "00000000";
                when "11011111" => rgb <= "00000000";
                when "11100000" => rgb <= "00000000";
                when "11100001" => rgb <= "00000000";
                when "11100010" => rgb <= "00000000";
                when "11100011" => rgb <= "00000000";
                when "11100100" => rgb <= "00000000";
                when "11100101" => rgb <= "00000000";
                when "11100110" => rgb <= "00000000";
                when "11100111" => rgb <= "00000000";
                when "11101000" => rgb <= "00000000";
                when "11101001" => rgb <= "00000000";
                when "11101010" => rgb <= "11101101";
                when "11101011" => rgb <= "11001111";
                when "11101100" => rgb <= "00000011";
                when "11101101" => rgb <= "00000000";
                when "11101110" => rgb <= "00000000";
                when "11101111" => rgb <= "00000010";
                when "11110000" => rgb <= "10111001";
                when "11110001" => rgb <= "11111110";
                when "11110010" => rgb <= "10101000";
                when "11110011" => rgb <= "00000000";
                when "11110100" => rgb <= "00000000";
                when "11110101" => rgb <= "00000000";
                when "11110110" => rgb <= "00000000";
                when "11110111" => rgb <= "00000000";
                when "11111000" => rgb <= "00000000";
                when "11111001" => rgb <= "00000000";
                when "11111010" => rgb <= "00000000";
                when "11111011" => rgb <= "00000000";
                when "11111100" => rgb <= "00000000";
                when "11111101" => rgb <= "00000000";
                when "11111110" => rgb <= "00000000";
                when "11111111" => rgb <= "00000000";
                when "100000000" => rgb <= "00000000";
                when "100000001" => rgb <= "00000000";
                when "100000010" => rgb <= "00000000";
                when "100000011" => rgb <= "00000000";
                when "100000100" => rgb <= "00000000";
                when "100000101" => rgb <= "00111001";
                when "100000110" => rgb <= "11111101";
                when "100000111" => rgb <= "10111011";
                when "100001000" => rgb <= "00000000";
                when "100001001" => rgb <= "00000000";
                when "100001010" => rgb <= "00000000";
                when "100001011" => rgb <= "00000000";
                when "100001100" => rgb <= "00110001";
                when "100001101" => rgb <= "11111110";
                when "100001110" => rgb <= "11111011";
                when "100001111" => rgb <= "01000011";
                when "100010000" => rgb <= "00000000";
                when "100010001" => rgb <= "00000000";
                when "100010010" => rgb <= "00000000";
                when "100010011" => rgb <= "00000000";
                when "100010100" => rgb <= "00000000";
                when "100010101" => rgb <= "00000000";
                when "100010110" => rgb <= "00000000";
                when "100010111" => rgb <= "00000000";
                when "100011000" => rgb <= "00000000";
                when "100011001" => rgb <= "00000000";
                when "100011010" => rgb <= "00000000";
                when "100011011" => rgb <= "00000000";
                when "100011100" => rgb <= "00000000";
                when "100011101" => rgb <= "00000000";
                when "100011110" => rgb <= "00000000";
                when "100011111" => rgb <= "00000000";
                when "100100000" => rgb <= "00000000";
                when "100100001" => rgb <= "10100011";
                when "100100010" => rgb <= "11111110";
                when "100100011" => rgb <= "01111010";
                when "100100100" => rgb <= "00000000";
                when "100100101" => rgb <= "00000000";
                when "100100110" => rgb <= "00000000";
                when "100100111" => rgb <= "00000000";
                when "100101000" => rgb <= "00001001";
                when "100101001" => rgb <= "10011101";
                when "100101010" => rgb <= "11111110";
                when "100101011" => rgb <= "10010110";
                when "100101100" => rgb <= "00000000";
                when "100101101" => rgb <= "00000000";
                when "100101110" => rgb <= "00000000";
                when "100101111" => rgb <= "00000000";
                when "100110000" => rgb <= "00000000";
                when "100110001" => rgb <= "00000000";
                when "100110010" => rgb <= "00000000";
                when "100110011" => rgb <= "00000000";
                when "100110100" => rgb <= "00000000";
                when "100110101" => rgb <= "00000000";
                when "100110110" => rgb <= "00000000";
                when "100110111" => rgb <= "00000000";
                when "100111000" => rgb <= "00000000";
                when "100111001" => rgb <= "00000000";
                when "100111010" => rgb <= "00000000";
                when "100111011" => rgb <= "00000000";
                when "100111100" => rgb <= "00000000";
                when "100111101" => rgb <= "11000110";
                when "100111110" => rgb <= "11110110";
                when "100111111" => rgb <= "00110110";
                when "101000000" => rgb <= "00000000";
                when "101000001" => rgb <= "00000000";
                when "101000010" => rgb <= "00000000";
                when "101000011" => rgb <= "00000000";
                when "101000100" => rgb <= "00000000";
                when "101000101" => rgb <= "00011110";
                when "101000110" => rgb <= "11100111";
                when "101000111" => rgb <= "11110110";
                when "101001000" => rgb <= "00100101";
                when "101001001" => rgb <= "00000000";
                when "101001010" => rgb <= "00000000";
                when "101001011" => rgb <= "00000000";
                when "101001100" => rgb <= "00000000";
                when "101001101" => rgb <= "00000000";
                when "101001110" => rgb <= "00000000";
                when "101001111" => rgb <= "00000000";
                when "101010000" => rgb <= "00000000";
                when "101010001" => rgb <= "00000000";
                when "101010010" => rgb <= "00000000";
                when "101010011" => rgb <= "00000000";
                when "101010100" => rgb <= "00000000";
                when "101010101" => rgb <= "00000000";
                when "101010110" => rgb <= "00000000";
                when "101010111" => rgb <= "00000000";
                when "101011000" => rgb <= "00000000";
                when "101011001" => rgb <= "11000110";
                when "101011010" => rgb <= "11101001";
                when "101011011" => rgb <= "00000000";
                when "101011100" => rgb <= "00000000";
                when "101011101" => rgb <= "00000000";
                when "101011110" => rgb <= "00000000";
                when "101011111" => rgb <= "00000000";
                when "101100000" => rgb <= "00000000";
                when "101100001" => rgb <= "00000000";
                when "101100010" => rgb <= "10011010";
                when "101100011" => rgb <= "11111110";
                when "101100100" => rgb <= "01001001";
                when "101100101" => rgb <= "00000000";
                when "101100110" => rgb <= "00000000";
                when "101100111" => rgb <= "00000000";
                when "101101000" => rgb <= "00000000";
                when "101101001" => rgb <= "00000000";
                when "101101010" => rgb <= "00000000";
                when "101101011" => rgb <= "00000000";
                when "101101100" => rgb <= "00000000";
                when "101101101" => rgb <= "00000000";
                when "101101110" => rgb <= "00000000";
                when "101101111" => rgb <= "00000000";
                when "101110000" => rgb <= "00000000";
                when "101110001" => rgb <= "00000000";
                when "101110010" => rgb <= "00000000";
                when "101110011" => rgb <= "00000000";
                when "101110100" => rgb <= "00001111";
                when "101110101" => rgb <= "11111110";
                when "101110110" => rgb <= "11101001";
                when "101110111" => rgb <= "00000000";
                when "101111000" => rgb <= "00000000";
                when "101111001" => rgb <= "00000000";
                when "101111010" => rgb <= "00000000";
                when "101111011" => rgb <= "00000000";
                when "101111100" => rgb <= "00000000";
                when "101111101" => rgb <= "00000000";
                when "101111110" => rgb <= "01111011";
                when "101111111" => rgb <= "11111110";
                when "110000000" => rgb <= "10000111";
                when "110000001" => rgb <= "00000000";
                when "110000010" => rgb <= "00000000";
                when "110000011" => rgb <= "00000000";
                when "110000100" => rgb <= "00000000";
                when "110000101" => rgb <= "00000000";
                when "110000110" => rgb <= "00000000";
                when "110000111" => rgb <= "00000000";
                when "110001000" => rgb <= "00000000";
                when "110001001" => rgb <= "00000000";
                when "110001010" => rgb <= "00000000";
                when "110001011" => rgb <= "00000000";
                when "110001100" => rgb <= "00000000";
                when "110001101" => rgb <= "00000000";
                when "110001110" => rgb <= "00000000";
                when "110001111" => rgb <= "00000000";
                when "110010000" => rgb <= "00001111";
                when "110010001" => rgb <= "11111110";
                when "110010010" => rgb <= "11101001";
                when "110010011" => rgb <= "00000000";
                when "110010100" => rgb <= "00000000";
                when "110010101" => rgb <= "00000000";
                when "110010110" => rgb <= "00000000";
                when "110010111" => rgb <= "00000000";
                when "110011000" => rgb <= "00000000";
                when "110011001" => rgb <= "00000000";
                when "110011010" => rgb <= "01111011";
                when "110011011" => rgb <= "11111110";
                when "110011100" => rgb <= "11000101";
                when "110011101" => rgb <= "00000000";
                when "110011110" => rgb <= "00000000";
                when "110011111" => rgb <= "00000000";
                when "110100000" => rgb <= "00000000";
                when "110100001" => rgb <= "00000000";
                when "110100010" => rgb <= "00000000";
                when "110100011" => rgb <= "00000000";
                when "110100100" => rgb <= "00000000";
                when "110100101" => rgb <= "00000000";
                when "110100110" => rgb <= "00000000";
                when "110100111" => rgb <= "00000000";
                when "110101000" => rgb <= "00000000";
                when "110101001" => rgb <= "00000000";
                when "110101010" => rgb <= "00000000";
                when "110101011" => rgb <= "00000000";
                when "110101100" => rgb <= "00001111";
                when "110101101" => rgb <= "11111110";
                when "110101110" => rgb <= "11001000";
                when "110101111" => rgb <= "00000000";
                when "110110000" => rgb <= "00000000";
                when "110110001" => rgb <= "00000000";
                when "110110010" => rgb <= "00000000";
                when "110110011" => rgb <= "00000000";
                when "110110100" => rgb <= "00000000";
                when "110110101" => rgb <= "00000000";
                when "110110110" => rgb <= "01000110";
                when "110110111" => rgb <= "11111110";
                when "110111000" => rgb <= "11100101";
                when "110111001" => rgb <= "00001000";
                when "110111010" => rgb <= "00000000";
                when "110111011" => rgb <= "00000000";
                when "110111100" => rgb <= "00000000";
                when "110111101" => rgb <= "00000000";
                when "110111110" => rgb <= "00000000";
                when "110111111" => rgb <= "00000000";
                when "111000000" => rgb <= "00000000";
                when "111000001" => rgb <= "00000000";
                when "111000010" => rgb <= "00000000";
                when "111000011" => rgb <= "00000000";
                when "111000100" => rgb <= "00000000";
                when "111000101" => rgb <= "00000000";
                when "111000110" => rgb <= "00000000";
                when "111000111" => rgb <= "00000000";
                when "111001000" => rgb <= "00001111";
                when "111001001" => rgb <= "11111110";
                when "111001010" => rgb <= "10100001";
                when "111001011" => rgb <= "00000000";
                when "111001100" => rgb <= "00000000";
                when "111001101" => rgb <= "00000000";
                when "111001110" => rgb <= "00000000";
                when "111001111" => rgb <= "00000000";
                when "111010000" => rgb <= "00000000";
                when "111010001" => rgb <= "00000000";
                when "111010010" => rgb <= "00110011";
                when "111010011" => rgb <= "11111110";
                when "111010100" => rgb <= "11111000";
                when "111010101" => rgb <= "00001101";
                when "111010110" => rgb <= "00000000";
                when "111010111" => rgb <= "00000000";
                when "111011000" => rgb <= "00000000";
                when "111011001" => rgb <= "00000000";
                when "111011010" => rgb <= "00000000";
                when "111011011" => rgb <= "00000000";
                when "111011100" => rgb <= "00000000";
                when "111011101" => rgb <= "00000000";
                when "111011110" => rgb <= "00000000";
                when "111011111" => rgb <= "00000000";
                when "111100000" => rgb <= "00000000";
                when "111100001" => rgb <= "00000000";
                when "111100010" => rgb <= "00000000";
                when "111100011" => rgb <= "00000000";
                when "111100100" => rgb <= "00001111";
                when "111100101" => rgb <= "11111110";
                when "111100110" => rgb <= "10100001";
                when "111100111" => rgb <= "00000000";
                when "111101000" => rgb <= "00000000";
                when "111101001" => rgb <= "00000000";
                when "111101010" => rgb <= "00000000";
                when "111101011" => rgb <= "00000000";
                when "111101100" => rgb <= "00000000";
                when "111101101" => rgb <= "00000000";
                when "111101110" => rgb <= "00110011";
                when "111101111" => rgb <= "11111110";
                when "111110000" => rgb <= "11111110";
                when "111110001" => rgb <= "00001110";
                when "111110010" => rgb <= "00000000";
                when "111110011" => rgb <= "00000000";
                when "111110100" => rgb <= "00000000";
                when "111110101" => rgb <= "00000000";
                when "111110110" => rgb <= "00000000";
                when "111110111" => rgb <= "00000000";
                when "111111000" => rgb <= "00000000";
                when "111111001" => rgb <= "00000000";
                when "111111010" => rgb <= "00000000";
                when "111111011" => rgb <= "00000000";
                when "111111100" => rgb <= "00000000";
                when "111111101" => rgb <= "00000000";
                when "111111110" => rgb <= "00000000";
                when "111111111" => rgb <= "00000000";
                when "1000000000" => rgb <= "00001010";
                when "1000000001" => rgb <= "11101010";
                when "1000000010" => rgb <= "10111010";
                when "1000000011" => rgb <= "00000000";
                when "1000000100" => rgb <= "00000000";
                when "1000000101" => rgb <= "00000000";
                when "1000000110" => rgb <= "00000000";
                when "1000000111" => rgb <= "00000000";
                when "1000001000" => rgb <= "00000000";
                when "1000001001" => rgb <= "00000000";
                when "1000001010" => rgb <= "01100001";
                when "1000001011" => rgb <= "11111110";
                when "1000001100" => rgb <= "11011010";
                when "1000001101" => rgb <= "00000101";
                when "1000001110" => rgb <= "00000000";
                when "1000001111" => rgb <= "00000000";
                when "1000010000" => rgb <= "00000000";
                when "1000010001" => rgb <= "00000000";
                when "1000010010" => rgb <= "00000000";
                when "1000010011" => rgb <= "00000000";
                when "1000010100" => rgb <= "00000000";
                when "1000010101" => rgb <= "00000000";
                when "1000010110" => rgb <= "00000000";
                when "1000010111" => rgb <= "00000000";
                when "1000011000" => rgb <= "00000000";
                when "1000011001" => rgb <= "00000000";
                when "1000011010" => rgb <= "00000000";
                when "1000011011" => rgb <= "00000000";
                when "1000011100" => rgb <= "00000000";
                when "1000011101" => rgb <= "11000110";
                when "1000011110" => rgb <= "11101110";
                when "1000011111" => rgb <= "00001100";
                when "1000100000" => rgb <= "00000000";
                when "1000100001" => rgb <= "00000000";
                when "1000100010" => rgb <= "00000000";
                when "1000100011" => rgb <= "00000000";
                when "1000100100" => rgb <= "00000000";
                when "1000100101" => rgb <= "00000011";
                when "1000100110" => rgb <= "10101100";
                when "1000100111" => rgb <= "11111110";
                when "1000101000" => rgb <= "10100000";
                when "1000101001" => rgb <= "00000000";
                when "1000101010" => rgb <= "00000000";
                when "1000101011" => rgb <= "00000000";
                when "1000101100" => rgb <= "00000000";
                when "1000101101" => rgb <= "00000000";
                when "1000101110" => rgb <= "00000000";
                when "1000101111" => rgb <= "00000000";
                when "1000110000" => rgb <= "00000000";
                when "1000110001" => rgb <= "00000000";
                when "1000110010" => rgb <= "00000000";
                when "1000110011" => rgb <= "00000000";
                when "1000110100" => rgb <= "00000000";
                when "1000110101" => rgb <= "00000000";
                when "1000110110" => rgb <= "00000000";
                when "1000110111" => rgb <= "00000000";
                when "1000111000" => rgb <= "00000000";
                when "1000111001" => rgb <= "01111011";
                when "1000111010" => rgb <= "11111110";
                when "1000111011" => rgb <= "10000011";
                when "1000111100" => rgb <= "00000001";
                when "1000111101" => rgb <= "00000000";
                when "1000111110" => rgb <= "00000000";
                when "1000111111" => rgb <= "00000000";
                when "1001000000" => rgb <= "00001100";
                when "1001000001" => rgb <= "10011101";
                when "1001000010" => rgb <= "11111110";
                when "1001000011" => rgb <= "11111000";
                when "1001000100" => rgb <= "00100101";
                when "1001000101" => rgb <= "00000000";
                when "1001000110" => rgb <= "00000000";
                when "1001000111" => rgb <= "00000000";
                when "1001001000" => rgb <= "00000000";
                when "1001001001" => rgb <= "00000000";
                when "1001001010" => rgb <= "00000000";
                when "1001001011" => rgb <= "00000000";
                when "1001001100" => rgb <= "00000000";
                when "1001001101" => rgb <= "00000000";
                when "1001001110" => rgb <= "00000000";
                when "1001001111" => rgb <= "00000000";
                when "1001010000" => rgb <= "00000000";
                when "1001010001" => rgb <= "00000000";
                when "1001010010" => rgb <= "00000000";
                when "1001010011" => rgb <= "00000000";
                when "1001010100" => rgb <= "00000000";
                when "1001010101" => rgb <= "00001010";
                when "1001010110" => rgb <= "11110000";
                when "1001010111" => rgb <= "100000000";
                when "1001011000" => rgb <= "10110110";
                when "1001011001" => rgb <= "01001101";
                when "1001011010" => rgb <= "01000001";
                when "1001011011" => rgb <= "10000000";
                when "1001011100" => rgb <= "11100101";
                when "1001011101" => rgb <= "100000000";
                when "1001011110" => rgb <= "11111110";
                when "1001011111" => rgb <= "01111010";
                when "1001100000" => rgb <= "00000000";
                when "1001100001" => rgb <= "00000000";
                when "1001100010" => rgb <= "00000000";
                when "1001100011" => rgb <= "00000000";
                when "1001100100" => rgb <= "00000000";
                when "1001100101" => rgb <= "00000000";
                when "1001100110" => rgb <= "00000000";
                when "1001100111" => rgb <= "00000000";
                when "1001101000" => rgb <= "00000000";
                when "1001101001" => rgb <= "00000000";
                when "1001101010" => rgb <= "00000000";
                when "1001101011" => rgb <= "00000000";
                when "1001101100" => rgb <= "00000000";
                when "1001101101" => rgb <= "00000000";
                when "1001101110" => rgb <= "00000000";
                when "1001101111" => rgb <= "00000000";
                when "1001110000" => rgb <= "00000000";
                when "1001110001" => rgb <= "00000000";
                when "1001110010" => rgb <= "00100111";
                when "1001110011" => rgb <= "11011000";
                when "1001110100" => rgb <= "11111110";
                when "1001110101" => rgb <= "11111110";
                when "1001110110" => rgb <= "11111110";
                when "1001110111" => rgb <= "11111110";
                when "1001111000" => rgb <= "11111110";
                when "1001111001" => rgb <= "11110001";
                when "1001111010" => rgb <= "01100110";
                when "1001111011" => rgb <= "00000001";
                when "1001111100" => rgb <= "00000000";
                when "1001111101" => rgb <= "00000000";
                when "1001111110" => rgb <= "00000000";
                when "1001111111" => rgb <= "00000000";
                when "1010000000" => rgb <= "00000000";
                when "1010000001" => rgb <= "00000000";
                when "1010000010" => rgb <= "00000000";
                when "1010000011" => rgb <= "00000000";
                when "1010000100" => rgb <= "00000000";
                when "1010000101" => rgb <= "00000000";
                when "1010000110" => rgb <= "00000000";
                when "1010000111" => rgb <= "00000000";
                when "1010001000" => rgb <= "00000000";
                when "1010001001" => rgb <= "00000000";
                when "1010001010" => rgb <= "00000000";
                when "1010001011" => rgb <= "00000000";
                when "1010001100" => rgb <= "00000000";
                when "1010001101" => rgb <= "00000000";
                when "1010001110" => rgb <= "00000000";
                when "1010001111" => rgb <= "00001010";
                when "1010010000" => rgb <= "10011100";
                when "1010010001" => rgb <= "11011110";
                when "1010010010" => rgb <= "11111110";
                when "1010010011" => rgb <= "11101001";
                when "1010010100" => rgb <= "10010110";
                when "1010010101" => rgb <= "00100011";
                when "1010010110" => rgb <= "00000000";
                when "1010010111" => rgb <= "00000000";
                when "1010011000" => rgb <= "00000000";
                when "1010011001" => rgb <= "00000000";
                when "1010011010" => rgb <= "00000000";
                when "1010011011" => rgb <= "00000000";
                when "1010011100" => rgb <= "00000000";
                when "1010011101" => rgb <= "00000000";
                when "1010011110" => rgb <= "00000000";
                when "1010011111" => rgb <= "00000000";
                when "1010100000" => rgb <= "00000000";
                when "1010100001" => rgb <= "00000000";
                when "1010100010" => rgb <= "00000000";
                when "1010100011" => rgb <= "00000000";
                when "1010100100" => rgb <= "00000000";
                when "1010100101" => rgb <= "00000000";
                when "1010100110" => rgb <= "00000000";
                when "1010100111" => rgb <= "00000000";
                when "1010101000" => rgb <= "00000000";
                when "1010101001" => rgb <= "00000000";
                when "1010101010" => rgb <= "00000000";
                when "1010101011" => rgb <= "00000000";
                when "1010101100" => rgb <= "00000000";
                when "1010101101" => rgb <= "00000000";
                when "1010101110" => rgb <= "00000000";
                when "1010101111" => rgb <= "00000000";
                when "1010110000" => rgb <= "00000000";
                when "1010110001" => rgb <= "00000000";
                when "1010110010" => rgb <= "00000000";
                when "1010110011" => rgb <= "00000000";
                when "1010110100" => rgb <= "00000000";
                when "1010110101" => rgb <= "00000000";
                when "1010110110" => rgb <= "00000000";
                when "1010110111" => rgb <= "00000000";
                when "1010111000" => rgb <= "00000000";
                when "1010111001" => rgb <= "00000000";
                when "1010111010" => rgb <= "00000000";
                when "1010111011" => rgb <= "00000000";
                when "1010111100" => rgb <= "00000000";
                when "1010111101" => rgb <= "00000000";
                when "1010111110" => rgb <= "00000000";
                when "1010111111" => rgb <= "00000000";
                when "1011000000" => rgb <= "00000000";
                when "1011000001" => rgb <= "00000000";
                when "1011000010" => rgb <= "00000000";
                when "1011000011" => rgb <= "00000000";
                when "1011000100" => rgb <= "00000000";
                when "1011000101" => rgb <= "00000000";
                when "1011000110" => rgb <= "00000000";
                when "1011000111" => rgb <= "00000000";
                when "1011001000" => rgb <= "00000000";
                when "1011001001" => rgb <= "00000000";
                when "1011001010" => rgb <= "00000000";
                when "1011001011" => rgb <= "00000000";
                when "1011001100" => rgb <= "00000000";
                when "1011001101" => rgb <= "00000000";
                when "1011001110" => rgb <= "00000000";
                when "1011001111" => rgb <= "00000000";
                when "1011010000" => rgb <= "00000000";
                when "1011010001" => rgb <= "00000000";
                when "1011010010" => rgb <= "00000000";
                when "1011010011" => rgb <= "00000000";
                when "1011010100" => rgb <= "00000000";
                when "1011010101" => rgb <= "00000000";
                when "1011010110" => rgb <= "00000000";
                when "1011010111" => rgb <= "00000000";
                when "1011011000" => rgb <= "00000000";
                when "1011011001" => rgb <= "00000000";
                when "1011011010" => rgb <= "00000000";
                when "1011011011" => rgb <= "00000000";
                when "1011011100" => rgb <= "00000000";
                when "1011011101" => rgb <= "00000000";
                when "1011011110" => rgb <= "00000000";
                when "1011011111" => rgb <= "00000000";
                when "1011100000" => rgb <= "00000000";
                when "1011100001" => rgb <= "00000000";
                when "1011100010" => rgb <= "00000000";
                when "1011100011" => rgb <= "00000000";
                when "1011100100" => rgb <= "00000000";
                when "1011100101" => rgb <= "00000000";
                when "1011100110" => rgb <= "00000000";
                when "1011100111" => rgb <= "00000000";
                when "1011101000" => rgb <= "00000000";
                when "1011101001" => rgb <= "00000000";
                when "1011101010" => rgb <= "00000000";
                when "1011101011" => rgb <= "00000000";
                when "1011101100" => rgb <= "00000000";
                when "1011101101" => rgb <= "00000000";
                when "1011101110" => rgb <= "00000000";
                when "1011101111" => rgb <= "00000000";
                when "1011110000" => rgb <= "00000000";
                when "1011110001" => rgb <= "00000000";
                when "1011110010" => rgb <= "00000000";
                when "1011110011" => rgb <= "00000000";
                when "1011110100" => rgb <= "00000000";
                when "1011110101" => rgb <= "00000000";
                when "1011110110" => rgb <= "00000000";
                when "1011110111" => rgb <= "00000000";
                when "1011111000" => rgb <= "00000000";
                when "1011111001" => rgb <= "00000000";
                when "1011111010" => rgb <= "00000000";
                when "1011111011" => rgb <= "00000000";
                when "1011111100" => rgb <= "00000000";
                when "1011111101" => rgb <= "00000000";
                when "1011111110" => rgb <= "00000000";
                when "1011111111" => rgb <= "00000000";
                when "1100000000" => rgb <= "00000000";
                when "1100000001" => rgb <= "00000000";
                when "1100000010" => rgb <= "00000000";
                when "1100000011" => rgb <= "00000000";
                when "1100000100" => rgb <= "00000000";
                when "1100000101" => rgb <= "00000000";
                when "1100000110" => rgb <= "00000000";
                when "1100000111" => rgb <= "00000000";
                when "1100001000" => rgb <= "00000000";
                when "1100001001" => rgb <= "00000000";
                when "1100001010" => rgb <= "00000000";
                when "1100001011" => rgb <= "00000000";
                when "1100001100" => rgb <= "00000000";
                when "1100001101" => rgb <= "00000000";
                when "1100001110" => rgb <= "00000000";
                when "1100001111" => rgb <= "00000000";
                when others => rgb <= "111111";
        end case;
    end if;
    end process;
    totaladr <= std_logic_vector(yadr) & std_logic_vector(xadr);
end;
