module weight_mem
    (
        input wire clk, 
        input wire reset,
        input wire [15:0] input_addr,
        output reg signed [7:0] weight_val
    );

    // 2^16 (size of neuron address) requires 65536 addresses
    reg signed [7:0] weight_mem[0:65535];

    // initializing input layer
    initial begin
        // layer 1 neuron 0
        weight_mem[16'h0000] <= 1;
        weight_mem[16'h0001] <= 0;
        weight_mem[16'h0002] <= 0;
        weight_mem[16'h0003] <= 0;
        weight_mem[16'h0004] <= 0;
        weight_mem[16'h0005] <= 0;
        weight_mem[16'h0006] <= 0;
        weight_mem[16'h0007] <= 0;
        weight_mem[16'h0008] <= 0;
        weight_mem[16'h0009] <= 0;
        weight_mem[16'h000A] <= 0;
        weight_mem[16'h000B] <= 0;
        weight_mem[16'h000C] <= 0;
        weight_mem[16'h000D] <= 0;
        weight_mem[16'h000E] <= 0;
        weight_mem[16'h000F] <= 0;
        weight_mem[16'h0010] <= 0;
        weight_mem[16'h0011] <= 0;
        weight_mem[16'h0012] <= 0;
        weight_mem[16'h0013] <= 0;
        weight_mem[16'h0014] <= 0;
        weight_mem[16'h0015] <= 0;
        weight_mem[16'h0016] <= 0;
        weight_mem[16'h0017] <= 0;
        weight_mem[16'h0018] <= 0;
        weight_mem[16'h0019] <= 0;
        weight_mem[16'h001A] <= 0;
        weight_mem[16'h001B] <= 0;
        weight_mem[16'h001C] <= 0;
        weight_mem[16'h001D] <= 0;
        weight_mem[16'h001E] <= 0;
        weight_mem[16'h001F] <= 0;
        weight_mem[16'h0020] <= 0;
        weight_mem[16'h0021] <= 0;
        weight_mem[16'h0022] <= 0;
        weight_mem[16'h0023] <= 0;
        weight_mem[16'h0024] <= 0;
        weight_mem[16'h0025] <= 0;
        weight_mem[16'h0026] <= 0;
        weight_mem[16'h0027] <= 0;
        weight_mem[16'h0028] <= 0;
        weight_mem[16'h0029] <= 0;
        weight_mem[16'h002A] <= 0;
        weight_mem[16'h002B] <= 0;
        weight_mem[16'h002C] <= 0;
        weight_mem[16'h002D] <= 0;
        weight_mem[16'h002E] <= 0;
        weight_mem[16'h002F] <= 0;
        weight_mem[16'h0030] <= 0;
        weight_mem[16'h0031] <= 0;
        weight_mem[16'h0032] <= 0;
        weight_mem[16'h0033] <= 0;
        weight_mem[16'h0034] <= 0;
        weight_mem[16'h0035] <= 0;
        weight_mem[16'h0036] <= 0;
        weight_mem[16'h0037] <= 0;
        weight_mem[16'h0038] <= 0;
        weight_mem[16'h0039] <= 0;
        weight_mem[16'h003A] <= 0;
        weight_mem[16'h003B] <= 0;
        weight_mem[16'h003C] <= 0;
        weight_mem[16'h003D] <= 0;
        weight_mem[16'h003E] <= 0;
        weight_mem[16'h003F] <= 0;
        weight_mem[16'h0040] <= 0;
        weight_mem[16'h0041] <= 0;
        weight_mem[16'h0042] <= 0;
        weight_mem[16'h0043] <= 0;
        weight_mem[16'h0044] <= 0;
        weight_mem[16'h0045] <= 0;
        weight_mem[16'h0046] <= 0;
        weight_mem[16'h0047] <= 0;
        weight_mem[16'h0048] <= 0;
        weight_mem[16'h0049] <= 0;
        weight_mem[16'h004A] <= 0;
        weight_mem[16'h004B] <= 0;
        weight_mem[16'h004C] <= 0;
        weight_mem[16'h004D] <= 0;
        weight_mem[16'h004E] <= 0;
        weight_mem[16'h004F] <= 0;
        weight_mem[16'h0050] <= 0;
        weight_mem[16'h0051] <= 0;
        weight_mem[16'h0052] <= 0;
        weight_mem[16'h0053] <= 0;
        weight_mem[16'h0054] <= 0;
        weight_mem[16'h0055] <= 0;
        weight_mem[16'h0056] <= 0;
        weight_mem[16'h0057] <= 0;
        weight_mem[16'h0058] <= 0;
        weight_mem[16'h0059] <= 0;
        weight_mem[16'h005A] <= 0;
        weight_mem[16'h005B] <= 0;
        weight_mem[16'h005C] <= 0;
        weight_mem[16'h005D] <= 0;
        weight_mem[16'h005E] <= 0;
        weight_mem[16'h005F] <= 0;
        weight_mem[16'h0060] <= 0;
        weight_mem[16'h0061] <= 0;
        weight_mem[16'h0062] <= 0;
        weight_mem[16'h0063] <= 0;
        weight_mem[16'h0064] <= 0;
        weight_mem[16'h0065] <= 0;
        weight_mem[16'h0066] <= 0;
        weight_mem[16'h0067] <= 0;
        weight_mem[16'h0068] <= 0;
        weight_mem[16'h0069] <= 0;
        weight_mem[16'h006A] <= 0;
        weight_mem[16'h006B] <= 0;
        weight_mem[16'h006C] <= 0;
        weight_mem[16'h006D] <= 0;
        weight_mem[16'h006E] <= 0;
        weight_mem[16'h006F] <= 0;
        weight_mem[16'h0070] <= 0;
        weight_mem[16'h0071] <= 0;
        weight_mem[16'h0072] <= 0;
        weight_mem[16'h0073] <= 0;
        weight_mem[16'h0074] <= 0;
        weight_mem[16'h0075] <= 0;
        weight_mem[16'h0076] <= 0;
        weight_mem[16'h0077] <= 0;
        weight_mem[16'h0078] <= 0;
        weight_mem[16'h0079] <= 0;
        weight_mem[16'h007A] <= 0;
        weight_mem[16'h007B] <= 0;
        weight_mem[16'h007C] <= 0;
        weight_mem[16'h007D] <= 0;
        weight_mem[16'h007E] <= 0;
        weight_mem[16'h007F] <= 0;
        weight_mem[16'h0080] <= 0;
        weight_mem[16'h0081] <= 0;
        weight_mem[16'h0082] <= 0;
        weight_mem[16'h0083] <= 0;
        weight_mem[16'h0084] <= 0;
        weight_mem[16'h0085] <= 0;
        weight_mem[16'h0086] <= 0;
        weight_mem[16'h0087] <= 0;
        weight_mem[16'h0088] <= 0;
        weight_mem[16'h0089] <= 0;
        weight_mem[16'h008A] <= 0;
        weight_mem[16'h008B] <= 0;
        weight_mem[16'h008C] <= 0;
        weight_mem[16'h008D] <= 0;
        weight_mem[16'h008E] <= 0;
        weight_mem[16'h008F] <= 0;
        weight_mem[16'h0090] <= 0;
        weight_mem[16'h0091] <= 0;
        weight_mem[16'h0092] <= 0;
        weight_mem[16'h0093] <= 0;
        weight_mem[16'h0094] <= 0;
        weight_mem[16'h0095] <= 0;
        weight_mem[16'h0096] <= 0;
        weight_mem[16'h0097] <= 0;
        weight_mem[16'h0098] <= 0;
        weight_mem[16'h0099] <= 0;
        weight_mem[16'h009A] <= 0;
        weight_mem[16'h009B] <= 0;
        weight_mem[16'h009C] <= 0;
        weight_mem[16'h009D] <= 0;
        weight_mem[16'h009E] <= 0;
        weight_mem[16'h009F] <= 0;
        weight_mem[16'h00A0] <= 0;
        weight_mem[16'h00A1] <= 0;
        weight_mem[16'h00A2] <= 0;
        weight_mem[16'h00A3] <= 0;
        weight_mem[16'h00A4] <= 0;
        weight_mem[16'h00A5] <= 0;
        weight_mem[16'h00A6] <= 0;
        weight_mem[16'h00A7] <= 0;
        weight_mem[16'h00A8] <= 0;
        weight_mem[16'h00A9] <= 0;
        weight_mem[16'h00AA] <= 0;
        weight_mem[16'h00AB] <= 0;
        weight_mem[16'h00AC] <= 0;
        weight_mem[16'h00AD] <= 0;
        weight_mem[16'h00AE] <= 0;
        weight_mem[16'h00AF] <= 0;
        weight_mem[16'h00B0] <= 0;
        weight_mem[16'h00B1] <= 0;
        weight_mem[16'h00B2] <= 0;
        weight_mem[16'h00B3] <= 0;
        weight_mem[16'h00B4] <= 0;
        weight_mem[16'h00B5] <= 0;
        weight_mem[16'h00B6] <= 0;
        weight_mem[16'h00B7] <= 0;
        weight_mem[16'h00B8] <= 0;
        weight_mem[16'h00B9] <= 0;
        weight_mem[16'h00BA] <= 0;
        weight_mem[16'h00BB] <= 0;
        weight_mem[16'h00BC] <= 0;
        weight_mem[16'h00BD] <= 0;
        weight_mem[16'h00BE] <= 0;
        weight_mem[16'h00BF] <= 0;
        weight_mem[16'h00C0] <= 0;
        weight_mem[16'h00C1] <= 0;
        weight_mem[16'h00C2] <= 0;
        weight_mem[16'h00C3] <= 0;
        weight_mem[16'h00C4] <= 0;
        weight_mem[16'h00C5] <= 0;
        weight_mem[16'h00C6] <= 0;
        weight_mem[16'h00C7] <= 0;
        weight_mem[16'h00C8] <= 0;
        weight_mem[16'h00C9] <= 0;
        weight_mem[16'h00CA] <= 0;
        weight_mem[16'h00CB] <= 0;
        weight_mem[16'h00CC] <= 0;
        weight_mem[16'h00CD] <= 0;
        weight_mem[16'h00CE] <= 0;
        weight_mem[16'h00CF] <= 0;
        weight_mem[16'h00D0] <= 0;
        weight_mem[16'h00D1] <= 0;
        weight_mem[16'h00D2] <= 0;
        weight_mem[16'h00D3] <= 0;
        weight_mem[16'h00D4] <= 0;
        weight_mem[16'h00D5] <= 0;
        weight_mem[16'h00D6] <= 0;
        weight_mem[16'h00D7] <= 0;
        weight_mem[16'h00D8] <= 0;
        weight_mem[16'h00D9] <= 0;
        weight_mem[16'h00DA] <= 0;
        weight_mem[16'h00DB] <= 0;
        weight_mem[16'h00DC] <= 0;
        weight_mem[16'h00DD] <= 0;
        weight_mem[16'h00DE] <= 0;
        weight_mem[16'h00DF] <= 0;
        weight_mem[16'h00E0] <= 0;
        weight_mem[16'h00E1] <= 0;
        weight_mem[16'h00E2] <= 0;
        weight_mem[16'h00E3] <= 0;
        weight_mem[16'h00E4] <= 0;
        weight_mem[16'h00E5] <= 0;
        weight_mem[16'h00E6] <= 0;
        weight_mem[16'h00E7] <= 0;
        weight_mem[16'h00E8] <= 0;
        weight_mem[16'h00E9] <= 0;
        weight_mem[16'h00EA] <= 0;
        weight_mem[16'h00EB] <= 0;
        weight_mem[16'h00EC] <= 0;
        weight_mem[16'h00ED] <= 0;
        weight_mem[16'h00EE] <= 0;
        weight_mem[16'h00EF] <= 0;
        weight_mem[16'h00F0] <= 0;
        weight_mem[16'h00F1] <= 0;
        weight_mem[16'h00F2] <= 0;
        weight_mem[16'h00F3] <= 0;
        weight_mem[16'h00F4] <= 0;
        weight_mem[16'h00F5] <= 0;
        weight_mem[16'h00F6] <= 0;
        weight_mem[16'h00F7] <= 0;
        weight_mem[16'h00F8] <= 0;
        weight_mem[16'h00F9] <= 0;
        weight_mem[16'h00FA] <= 0;
        weight_mem[16'h00FB] <= 0;
        weight_mem[16'h00FC] <= 0;
        weight_mem[16'h00FD] <= 0;
        weight_mem[16'h00FE] <= 0;
        weight_mem[16'h00FF] <= 0;
        weight_mem[16'h0100] <= 0;
        weight_mem[16'h0101] <= 0;
        weight_mem[16'h0102] <= 0;
        weight_mem[16'h0103] <= 0;
        weight_mem[16'h0104] <= 0;
        weight_mem[16'h0105] <= 0;
        weight_mem[16'h0106] <= 0;
        weight_mem[16'h0107] <= 0;
        weight_mem[16'h0108] <= 0;
        weight_mem[16'h0109] <= 0;
        weight_mem[16'h010A] <= 0;
        weight_mem[16'h010B] <= 0;
        weight_mem[16'h010C] <= 0;
        weight_mem[16'h010D] <= 0;
        weight_mem[16'h010E] <= 0;
        weight_mem[16'h010F] <= 0;
        weight_mem[16'h0110] <= 0;
        weight_mem[16'h0111] <= 0;
        weight_mem[16'h0112] <= 0;
        weight_mem[16'h0113] <= 0;
        weight_mem[16'h0114] <= 0;
        weight_mem[16'h0115] <= 0;
        weight_mem[16'h0116] <= 0;
        weight_mem[16'h0117] <= 0;
        weight_mem[16'h0118] <= 0;
        weight_mem[16'h0119] <= 0;
        weight_mem[16'h011A] <= 0;
        weight_mem[16'h011B] <= 0;
        weight_mem[16'h011C] <= 0;
        weight_mem[16'h011D] <= 0;
        weight_mem[16'h011E] <= 0;
        weight_mem[16'h011F] <= 0;
        weight_mem[16'h0120] <= 0;
        weight_mem[16'h0121] <= 0;
        weight_mem[16'h0122] <= 0;
        weight_mem[16'h0123] <= 0;
        weight_mem[16'h0124] <= 0;
        weight_mem[16'h0125] <= 0;
        weight_mem[16'h0126] <= 0;
        weight_mem[16'h0127] <= 0;
        weight_mem[16'h0128] <= 0;
        weight_mem[16'h0129] <= 0;
        weight_mem[16'h012A] <= 0;
        weight_mem[16'h012B] <= 0;
        weight_mem[16'h012C] <= 0;
        weight_mem[16'h012D] <= 0;
        weight_mem[16'h012E] <= 0;
        weight_mem[16'h012F] <= 0;
        weight_mem[16'h0130] <= 0;
        weight_mem[16'h0131] <= 0;
        weight_mem[16'h0132] <= 0;
        weight_mem[16'h0133] <= 0;
        weight_mem[16'h0134] <= 0;
        weight_mem[16'h0135] <= 0;
        weight_mem[16'h0136] <= 0;
        weight_mem[16'h0137] <= 0;
        weight_mem[16'h0138] <= 0;
        weight_mem[16'h0139] <= 0;
        weight_mem[16'h013A] <= 0;
        weight_mem[16'h013B] <= 0;
        weight_mem[16'h013C] <= 0;
        weight_mem[16'h013D] <= 0;
        weight_mem[16'h013E] <= 0;
        weight_mem[16'h013F] <= 0;
        weight_mem[16'h0140] <= 0;
        weight_mem[16'h0141] <= 0;
        weight_mem[16'h0142] <= 0;
        weight_mem[16'h0143] <= 0;
        weight_mem[16'h0144] <= 0;
        weight_mem[16'h0145] <= 0;
        weight_mem[16'h0146] <= 0;
        weight_mem[16'h0147] <= 0;
        weight_mem[16'h0148] <= 0;
        weight_mem[16'h0149] <= 0;
        weight_mem[16'h014A] <= 0;
        weight_mem[16'h014B] <= 0;
        weight_mem[16'h014C] <= 0;
        weight_mem[16'h014D] <= 0;
        weight_mem[16'h014E] <= 0;
        weight_mem[16'h014F] <= 0;
        weight_mem[16'h0150] <= 0;
        weight_mem[16'h0151] <= 0;
        weight_mem[16'h0152] <= 0;
        weight_mem[16'h0153] <= 0;
        weight_mem[16'h0154] <= 0;
        weight_mem[16'h0155] <= 0;
        weight_mem[16'h0156] <= 0;
        weight_mem[16'h0157] <= 0;
        weight_mem[16'h0158] <= 0;
        weight_mem[16'h0159] <= 0;
        weight_mem[16'h015A] <= 0;
        weight_mem[16'h015B] <= 0;
        weight_mem[16'h015C] <= 0;
        weight_mem[16'h015D] <= 0;
        weight_mem[16'h015E] <= 0;
        weight_mem[16'h015F] <= 0;
        weight_mem[16'h0160] <= 0;
        weight_mem[16'h0161] <= 0;
        weight_mem[16'h0162] <= 0;
        weight_mem[16'h0163] <= 0;
        weight_mem[16'h0164] <= 0;
        weight_mem[16'h0165] <= 0;
        weight_mem[16'h0166] <= 0;
        weight_mem[16'h0167] <= 0;
        weight_mem[16'h0168] <= 0;
        weight_mem[16'h0169] <= 0;
        weight_mem[16'h016A] <= 0;
        weight_mem[16'h016B] <= 0;
        weight_mem[16'h016C] <= 0;
        weight_mem[16'h016D] <= 0;
        weight_mem[16'h016E] <= 0;
        weight_mem[16'h016F] <= 0;
        weight_mem[16'h0170] <= 0;
        weight_mem[16'h0171] <= 0;
        weight_mem[16'h0172] <= 0;
        weight_mem[16'h0173] <= 0;
        weight_mem[16'h0174] <= 0;
        weight_mem[16'h0175] <= 0;
        weight_mem[16'h0176] <= 0;
        weight_mem[16'h0177] <= 0;
        weight_mem[16'h0178] <= 0;
        weight_mem[16'h0179] <= 0;
        weight_mem[16'h017A] <= 0;
        weight_mem[16'h017B] <= 0;
        weight_mem[16'h017C] <= 0;
        weight_mem[16'h017D] <= 0;
        weight_mem[16'h017E] <= 0;
        weight_mem[16'h017F] <= 0;
        weight_mem[16'h0180] <= 0;
        weight_mem[16'h0181] <= 0;
        weight_mem[16'h0182] <= 0;
        weight_mem[16'h0183] <= 0;
        weight_mem[16'h0184] <= 0;
        weight_mem[16'h0185] <= 0;
        weight_mem[16'h0186] <= 0;
        weight_mem[16'h0187] <= 0;
        weight_mem[16'h0188] <= 0;
        weight_mem[16'h0189] <= 0;
        weight_mem[16'h018A] <= 0;
        weight_mem[16'h018B] <= 0;
        weight_mem[16'h018C] <= 0;
        weight_mem[16'h018D] <= 0;
        weight_mem[16'h018E] <= 0;
        weight_mem[16'h018F] <= 0;
        weight_mem[16'h0190] <= 0;
        weight_mem[16'h0191] <= 0;
        weight_mem[16'h0192] <= 0;
        weight_mem[16'h0193] <= 0;
        weight_mem[16'h0194] <= 0;
        weight_mem[16'h0195] <= 0;
        weight_mem[16'h0196] <= 0;
        weight_mem[16'h0197] <= 0;
        weight_mem[16'h0198] <= 0;
        weight_mem[16'h0199] <= 0;
        weight_mem[16'h019A] <= 0;
        weight_mem[16'h019B] <= 0;
        weight_mem[16'h019C] <= 0;
        weight_mem[16'h019D] <= 0;
        weight_mem[16'h019E] <= 0;
        weight_mem[16'h019F] <= 0;
        weight_mem[16'h01A0] <= 0;
        weight_mem[16'h01A1] <= 0;
        weight_mem[16'h01A2] <= 0;
        weight_mem[16'h01A3] <= 0;
        weight_mem[16'h01A4] <= 0;
        weight_mem[16'h01A5] <= 0;
        weight_mem[16'h01A6] <= 0;
        weight_mem[16'h01A7] <= 0;
        weight_mem[16'h01A8] <= 0;
        weight_mem[16'h01A9] <= 0;
        weight_mem[16'h01AA] <= 0;
        weight_mem[16'h01AB] <= 0;
        weight_mem[16'h01AC] <= 0;
        weight_mem[16'h01AD] <= 0;
        weight_mem[16'h01AE] <= 0;
        weight_mem[16'h01AF] <= 0;

        // layer 1 neuron 1
        weight_mem[16'h0200] <= 0;
        weight_mem[16'h0201] <= 0;
        weight_mem[16'h0202] <= 0;
        weight_mem[16'h0203] <= 0;
        weight_mem[16'h0204] <= 0;
        weight_mem[16'h0205] <= 0;
        weight_mem[16'h0206] <= 0;
        weight_mem[16'h0207] <= 0;
        weight_mem[16'h0208] <= 0;
        weight_mem[16'h0209] <= 0;
        weight_mem[16'h020A] <= 0;
        weight_mem[16'h020B] <= 0;
        weight_mem[16'h020C] <= 0;
        weight_mem[16'h020D] <= 0;
        weight_mem[16'h020E] <= 0;
        weight_mem[16'h020F] <= 0;
        weight_mem[16'h0210] <= 0;
        weight_mem[16'h0211] <= 0;
        weight_mem[16'h0212] <= 0;
        weight_mem[16'h0213] <= 0;
        weight_mem[16'h0214] <= 0;
        weight_mem[16'h0215] <= 0;
        weight_mem[16'h0216] <= 0;
        weight_mem[16'h0217] <= 0;
        weight_mem[16'h0218] <= 0;
        weight_mem[16'h0219] <= 0;
        weight_mem[16'h021A] <= 0;
        weight_mem[16'h021B] <= 0;
        weight_mem[16'h021C] <= 0;
        weight_mem[16'h021D] <= 0;
        weight_mem[16'h021E] <= 0;
        weight_mem[16'h021F] <= 0;
        weight_mem[16'h0220] <= 0;
        weight_mem[16'h0221] <= 0;
        weight_mem[16'h0222] <= 0;
        weight_mem[16'h0223] <= 0;
        weight_mem[16'h0224] <= 0;
        weight_mem[16'h0225] <= 0;
        weight_mem[16'h0226] <= 0;
        weight_mem[16'h0227] <= 0;
        weight_mem[16'h0228] <= 0;
        weight_mem[16'h0229] <= 0;
        weight_mem[16'h022A] <= 0;
        weight_mem[16'h022B] <= 0;
        weight_mem[16'h022C] <= 0;
        weight_mem[16'h022D] <= 0;
        weight_mem[16'h022E] <= 0;
        weight_mem[16'h022F] <= 0;
        weight_mem[16'h0230] <= 0;
        weight_mem[16'h0231] <= 0;
        weight_mem[16'h0232] <= 0;
        weight_mem[16'h0233] <= 0;
        weight_mem[16'h0234] <= 0;
        weight_mem[16'h0235] <= 0;
        weight_mem[16'h0236] <= 0;
        weight_mem[16'h0237] <= 0;
        weight_mem[16'h0238] <= 0;
        weight_mem[16'h0239] <= 0;
        weight_mem[16'h023A] <= 0;
        weight_mem[16'h023B] <= 0;
        weight_mem[16'h023C] <= 0;
        weight_mem[16'h023D] <= 0;
        weight_mem[16'h023E] <= 0;
        weight_mem[16'h023F] <= 0;
        weight_mem[16'h0240] <= 0;
        weight_mem[16'h0241] <= 0;
        weight_mem[16'h0242] <= 0;
        weight_mem[16'h0243] <= 0;
        weight_mem[16'h0244] <= 0;
        weight_mem[16'h0245] <= 0;
        weight_mem[16'h0246] <= 0;
        weight_mem[16'h0247] <= 0;
        weight_mem[16'h0248] <= 0;
        weight_mem[16'h0249] <= 0;
        weight_mem[16'h024A] <= 0;
        weight_mem[16'h024B] <= 0;
        weight_mem[16'h024C] <= 0;
        weight_mem[16'h024D] <= 0;
        weight_mem[16'h024E] <= 0;
        weight_mem[16'h024F] <= 0;
        weight_mem[16'h0250] <= 0;
        weight_mem[16'h0251] <= 0;
        weight_mem[16'h0252] <= 0;
        weight_mem[16'h0253] <= 0;
        weight_mem[16'h0254] <= 0;
        weight_mem[16'h0255] <= 0;
        weight_mem[16'h0256] <= 0;
        weight_mem[16'h0257] <= 0;
        weight_mem[16'h0258] <= 0;
        weight_mem[16'h0259] <= 0;
        weight_mem[16'h025A] <= 0;
        weight_mem[16'h025B] <= 0;
        weight_mem[16'h025C] <= 0;
        weight_mem[16'h025D] <= 0;
        weight_mem[16'h025E] <= 0;
        weight_mem[16'h025F] <= 0;
        weight_mem[16'h0260] <= 0;
        weight_mem[16'h0261] <= 0;
        weight_mem[16'h0262] <= 0;
        weight_mem[16'h0263] <= 0;
        weight_mem[16'h0264] <= 0;
        weight_mem[16'h0265] <= 0;
        weight_mem[16'h0266] <= 0;
        weight_mem[16'h0267] <= 0;
        weight_mem[16'h0268] <= 0;
        weight_mem[16'h0269] <= 0;
        weight_mem[16'h026A] <= 0;
        weight_mem[16'h026B] <= 0;
        weight_mem[16'h026C] <= 0;
        weight_mem[16'h026D] <= 0;
        weight_mem[16'h026E] <= 0;
        weight_mem[16'h026F] <= 0;
        weight_mem[16'h0270] <= 0;
        weight_mem[16'h0271] <= 0;
        weight_mem[16'h0272] <= 0;
        weight_mem[16'h0273] <= 0;
        weight_mem[16'h0274] <= 0;
        weight_mem[16'h0275] <= 0;
        weight_mem[16'h0276] <= 0;
        weight_mem[16'h0277] <= 0;
        weight_mem[16'h0278] <= 0;
        weight_mem[16'h0279] <= 0;
        weight_mem[16'h027A] <= 0;
        weight_mem[16'h027B] <= 0;
        weight_mem[16'h027C] <= 0;
        weight_mem[16'h027D] <= 0;
        weight_mem[16'h027E] <= 0;
        weight_mem[16'h027F] <= 0;
        weight_mem[16'h0280] <= 0;
        weight_mem[16'h0281] <= 0;
        weight_mem[16'h0282] <= 0;
        weight_mem[16'h0283] <= 0;
        weight_mem[16'h0284] <= 0;
        weight_mem[16'h0285] <= 0;
        weight_mem[16'h0286] <= 0;
        weight_mem[16'h0287] <= 0;
        weight_mem[16'h0288] <= 0;
        weight_mem[16'h0289] <= 0;
        weight_mem[16'h028A] <= 0;
        weight_mem[16'h028B] <= 0;
        weight_mem[16'h028C] <= 0;
        weight_mem[16'h028D] <= 0;
        weight_mem[16'h028E] <= 0;
        weight_mem[16'h028F] <= 0;
        weight_mem[16'h0290] <= 0;
        weight_mem[16'h0291] <= 0;
        weight_mem[16'h0292] <= 0;
        weight_mem[16'h0293] <= 0;
        weight_mem[16'h0294] <= 0;
        weight_mem[16'h0295] <= 0;
        weight_mem[16'h0296] <= 0;
        weight_mem[16'h0297] <= 0;
        weight_mem[16'h0298] <= 0;
        weight_mem[16'h0299] <= 0;
        weight_mem[16'h029A] <= 0;
        weight_mem[16'h029B] <= 0;
        weight_mem[16'h029C] <= 0;
        weight_mem[16'h029D] <= 0;
        weight_mem[16'h029E] <= 0;
        weight_mem[16'h029F] <= 0;
        weight_mem[16'h02A0] <= 0;
        weight_mem[16'h02A1] <= 0;
        weight_mem[16'h02A2] <= 0;
        weight_mem[16'h02A3] <= 0;
        weight_mem[16'h02A4] <= 0;
        weight_mem[16'h02A5] <= 0;
        weight_mem[16'h02A6] <= 0;
        weight_mem[16'h02A7] <= 0;
        weight_mem[16'h02A8] <= 0;
        weight_mem[16'h02A9] <= 0;
        weight_mem[16'h02AA] <= 0;
        weight_mem[16'h02AB] <= 0;
        weight_mem[16'h02AC] <= 0;
        weight_mem[16'h02AD] <= 0;
        weight_mem[16'h02AE] <= 0;
        weight_mem[16'h02AF] <= 0;
        weight_mem[16'h02B0] <= 0;
        weight_mem[16'h02B1] <= 0;
        weight_mem[16'h02B2] <= 0;
        weight_mem[16'h02B3] <= 0;
        weight_mem[16'h02B4] <= 0;
        weight_mem[16'h02B5] <= 0;
        weight_mem[16'h02B6] <= 0;
        weight_mem[16'h02B7] <= 0;
        weight_mem[16'h02B8] <= 0;
        weight_mem[16'h02B9] <= 0;
        weight_mem[16'h02BA] <= 0;
        weight_mem[16'h02BB] <= 0;
        weight_mem[16'h02BC] <= 0;
        weight_mem[16'h02BD] <= 0;
        weight_mem[16'h02BE] <= 0;
        weight_mem[16'h02BF] <= 0;
        weight_mem[16'h02C0] <= 0;
        weight_mem[16'h02C1] <= 0;
        weight_mem[16'h02C2] <= 0;
        weight_mem[16'h02C3] <= 0;
        weight_mem[16'h02C4] <= 0;
        weight_mem[16'h02C5] <= 0;
        weight_mem[16'h02C6] <= 0;
        weight_mem[16'h02C7] <= 0;
        weight_mem[16'h02C8] <= 0;
        weight_mem[16'h02C9] <= 0;
        weight_mem[16'h02CA] <= 0;
        weight_mem[16'h02CB] <= 0;
        weight_mem[16'h02CC] <= 0;
        weight_mem[16'h02CD] <= 0;
        weight_mem[16'h02CE] <= 0;
        weight_mem[16'h02CF] <= 0;
        weight_mem[16'h02D0] <= 0;
        weight_mem[16'h02D1] <= 0;
        weight_mem[16'h02D2] <= 0;
        weight_mem[16'h02D3] <= 0;
        weight_mem[16'h02D4] <= 0;
        weight_mem[16'h02D5] <= 0;
        weight_mem[16'h02D6] <= 0;
        weight_mem[16'h02D7] <= 0;
        weight_mem[16'h02D8] <= 0;
        weight_mem[16'h02D9] <= 0;
        weight_mem[16'h02DA] <= 0;
        weight_mem[16'h02DB] <= 0;
        weight_mem[16'h02DC] <= 0;
        weight_mem[16'h02DD] <= 0;
        weight_mem[16'h02DE] <= 0;
        weight_mem[16'h02DF] <= 0;
        weight_mem[16'h02E0] <= 0;
        weight_mem[16'h02E1] <= 0;
        weight_mem[16'h02E2] <= 0;
        weight_mem[16'h02E3] <= 0;
        weight_mem[16'h02E4] <= 0;
        weight_mem[16'h02E5] <= 0;
        weight_mem[16'h02E6] <= 0;
        weight_mem[16'h02E7] <= 0;
        weight_mem[16'h02E8] <= 0;
        weight_mem[16'h02E9] <= 0;
        weight_mem[16'h02EA] <= 0;
        weight_mem[16'h02EB] <= 0;
        weight_mem[16'h02EC] <= 0;
        weight_mem[16'h02ED] <= 0;
        weight_mem[16'h02EE] <= 0;
        weight_mem[16'h02EF] <= 0;
        weight_mem[16'h02F0] <= 0;
        weight_mem[16'h02F1] <= 0;
        weight_mem[16'h02F2] <= 0;
        weight_mem[16'h02F3] <= 0;
        weight_mem[16'h02F4] <= 0;
        weight_mem[16'h02F5] <= 0;
        weight_mem[16'h02F6] <= 0;
        weight_mem[16'h02F7] <= 0;
        weight_mem[16'h02F8] <= 0;
        weight_mem[16'h02F9] <= 0;
        weight_mem[16'h02FA] <= 0;
        weight_mem[16'h02FB] <= 0;
        weight_mem[16'h02FC] <= 0;
        weight_mem[16'h02FD] <= 0;
        weight_mem[16'h02FE] <= 0;
        weight_mem[16'h02FF] <= 0;
        weight_mem[16'h0300] <= 0;
        weight_mem[16'h0301] <= 0;
        weight_mem[16'h0302] <= 0;
        weight_mem[16'h0303] <= 0;
        weight_mem[16'h0304] <= 0;
        weight_mem[16'h0305] <= 0;
        weight_mem[16'h0306] <= 0;
        weight_mem[16'h0307] <= 0;
        weight_mem[16'h0308] <= 0;
        weight_mem[16'h0309] <= 0;
        weight_mem[16'h030A] <= 0;
        weight_mem[16'h030B] <= 0;
        weight_mem[16'h030C] <= 0;
        weight_mem[16'h030D] <= 0;
        weight_mem[16'h030E] <= 0;
        weight_mem[16'h030F] <= 0;
        weight_mem[16'h0310] <= 0;
        weight_mem[16'h0311] <= 0;
        weight_mem[16'h0312] <= 0;
        weight_mem[16'h0313] <= 0;
        weight_mem[16'h0314] <= 0;
        weight_mem[16'h0315] <= 0;
        weight_mem[16'h0316] <= 0;
        weight_mem[16'h0317] <= 0;
        weight_mem[16'h0318] <= 0;
        weight_mem[16'h0319] <= 0;
        weight_mem[16'h031A] <= 0;
        weight_mem[16'h031B] <= 0;
        weight_mem[16'h031C] <= 0;
        weight_mem[16'h031D] <= 0;
        weight_mem[16'h031E] <= 0;
        weight_mem[16'h031F] <= 0;
        weight_mem[16'h0320] <= 0;
        weight_mem[16'h0321] <= 0;
        weight_mem[16'h0322] <= 0;
        weight_mem[16'h0323] <= 0;
        weight_mem[16'h0324] <= 0;
        weight_mem[16'h0325] <= 0;
        weight_mem[16'h0326] <= 0;
        weight_mem[16'h0327] <= 0;
        weight_mem[16'h0328] <= 0;
        weight_mem[16'h0329] <= 0;
        weight_mem[16'h032A] <= 0;
        weight_mem[16'h032B] <= 0;
        weight_mem[16'h032C] <= 0;
        weight_mem[16'h032D] <= 0;
        weight_mem[16'h032E] <= 0;
        weight_mem[16'h032F] <= 0;
        weight_mem[16'h0330] <= 0;
        weight_mem[16'h0331] <= 0;
        weight_mem[16'h0332] <= 0;
        weight_mem[16'h0333] <= 0;
        weight_mem[16'h0334] <= 0;
        weight_mem[16'h0335] <= 0;
        weight_mem[16'h0336] <= 0;
        weight_mem[16'h0337] <= 0;
        weight_mem[16'h0338] <= 0;
        weight_mem[16'h0339] <= 0;
        weight_mem[16'h033A] <= 0;
        weight_mem[16'h033B] <= 0;
        weight_mem[16'h033C] <= 0;
        weight_mem[16'h033D] <= 0;
        weight_mem[16'h033E] <= 0;
        weight_mem[16'h033F] <= 0;
        weight_mem[16'h0340] <= 0;
        weight_mem[16'h0341] <= 0;
        weight_mem[16'h0342] <= 0;
        weight_mem[16'h0343] <= 0;
        weight_mem[16'h0344] <= 0;
        weight_mem[16'h0345] <= 0;
        weight_mem[16'h0346] <= 0;
        weight_mem[16'h0347] <= 0;
        weight_mem[16'h0348] <= 0;
        weight_mem[16'h0349] <= 0;
        weight_mem[16'h034A] <= 0;
        weight_mem[16'h034B] <= 0;
        weight_mem[16'h034C] <= 0;
        weight_mem[16'h034D] <= 0;
        weight_mem[16'h034E] <= 0;
        weight_mem[16'h034F] <= 0;
        weight_mem[16'h0350] <= 0;
        weight_mem[16'h0351] <= 0;
        weight_mem[16'h0352] <= 0;
        weight_mem[16'h0353] <= 0;
        weight_mem[16'h0354] <= 0;
        weight_mem[16'h0355] <= 0;
        weight_mem[16'h0356] <= 0;
        weight_mem[16'h0357] <= 0;
        weight_mem[16'h0358] <= 0;
        weight_mem[16'h0359] <= 0;
        weight_mem[16'h035A] <= 0;
        weight_mem[16'h035B] <= 0;
        weight_mem[16'h035C] <= 0;
        weight_mem[16'h035D] <= 0;
        weight_mem[16'h035E] <= 0;
        weight_mem[16'h035F] <= 0;
        weight_mem[16'h0360] <= 0;
        weight_mem[16'h0361] <= 0;
        weight_mem[16'h0362] <= 0;
        weight_mem[16'h0363] <= 0;
        weight_mem[16'h0364] <= 0;
        weight_mem[16'h0365] <= 0;
        weight_mem[16'h0366] <= 0;
        weight_mem[16'h0367] <= 0;
        weight_mem[16'h0368] <= 0;
        weight_mem[16'h0369] <= 0;
        weight_mem[16'h036A] <= 0;
        weight_mem[16'h036B] <= 0;
        weight_mem[16'h036C] <= 0;
        weight_mem[16'h036D] <= 0;
        weight_mem[16'h036E] <= 0;
        weight_mem[16'h036F] <= 0;
        weight_mem[16'h0370] <= 0;
        weight_mem[16'h0371] <= 0;
        weight_mem[16'h0372] <= 0;
        weight_mem[16'h0373] <= 0;
        weight_mem[16'h0374] <= 0;
        weight_mem[16'h0375] <= 0;
        weight_mem[16'h0376] <= 0;
        weight_mem[16'h0377] <= 0;
        weight_mem[16'h0378] <= 0;
        weight_mem[16'h0379] <= 0;
        weight_mem[16'h037A] <= 0;
        weight_mem[16'h037B] <= 0;
        weight_mem[16'h037C] <= 0;
        weight_mem[16'h037D] <= 0;
        weight_mem[16'h037E] <= 0;
        weight_mem[16'h037F] <= 0;
        weight_mem[16'h0380] <= 0;
        weight_mem[16'h0381] <= 0;
        weight_mem[16'h0382] <= 0;
        weight_mem[16'h0383] <= 0;
        weight_mem[16'h0384] <= 0;
        weight_mem[16'h0385] <= 0;
        weight_mem[16'h0386] <= 0;
        weight_mem[16'h0387] <= 0;
        weight_mem[16'h0388] <= 0;
        weight_mem[16'h0389] <= 0;
        weight_mem[16'h038A] <= 0;
        weight_mem[16'h038B] <= 0;
        weight_mem[16'h038C] <= 0;
        weight_mem[16'h038D] <= 0;
        weight_mem[16'h038E] <= 0;
        weight_mem[16'h038F] <= 0;
        weight_mem[16'h0390] <= 0;
        weight_mem[16'h0391] <= 0;
        weight_mem[16'h0392] <= 0;
        weight_mem[16'h0393] <= 0;
        weight_mem[16'h0394] <= 0;
        weight_mem[16'h0395] <= 0;
        weight_mem[16'h0396] <= 0;
        weight_mem[16'h0397] <= 0;
        weight_mem[16'h0398] <= 0;
        weight_mem[16'h0399] <= 0;
        weight_mem[16'h039A] <= 0;
        weight_mem[16'h039B] <= 0;
        weight_mem[16'h039C] <= 0;
        weight_mem[16'h039D] <= 0;
        weight_mem[16'h039E] <= 0;
        weight_mem[16'h039F] <= 0;
        weight_mem[16'h03A0] <= 0;
        weight_mem[16'h03A1] <= 0;
        weight_mem[16'h03A2] <= 0;
        weight_mem[16'h03A3] <= 0;
        weight_mem[16'h03A4] <= 0;
        weight_mem[16'h03A5] <= 0;
        weight_mem[16'h03A6] <= 0;
        weight_mem[16'h03A7] <= 0;
        weight_mem[16'h03A8] <= 0;
        weight_mem[16'h03A9] <= 0;
        weight_mem[16'h03AA] <= 0;
        weight_mem[16'h03AB] <= 0;
        weight_mem[16'h03AC] <= 0;
        weight_mem[16'h03AD] <= 0;
        weight_mem[16'h03AE] <= 0;
        weight_mem[16'h03AF] <= 0;

        // layer 1 neuron 2
        weight_mem[16'h0400] <= 0;
        weight_mem[16'h0401] <= 0;
        weight_mem[16'h0402] <= 0;
        weight_mem[16'h0403] <= 0;
        weight_mem[16'h0404] <= 0;
        weight_mem[16'h0405] <= 0;
        weight_mem[16'h0406] <= 0;
        weight_mem[16'h0407] <= 0;
        weight_mem[16'h0408] <= 0;
        weight_mem[16'h0409] <= 0;
        weight_mem[16'h040A] <= 0;
        weight_mem[16'h040B] <= 0;
        weight_mem[16'h040C] <= 0;
        weight_mem[16'h040D] <= 0;
        weight_mem[16'h040E] <= 0;
        weight_mem[16'h040F] <= 0;
        weight_mem[16'h0410] <= 0;
        weight_mem[16'h0411] <= 0;
        weight_mem[16'h0412] <= 0;
        weight_mem[16'h0413] <= 0;
        weight_mem[16'h0414] <= 0;
        weight_mem[16'h0415] <= 0;
        weight_mem[16'h0416] <= 0;
        weight_mem[16'h0417] <= 0;
        weight_mem[16'h0418] <= 0;
        weight_mem[16'h0419] <= 0;
        weight_mem[16'h041A] <= 0;
        weight_mem[16'h041B] <= 0;
        weight_mem[16'h041C] <= 0;
        weight_mem[16'h041D] <= 0;
        weight_mem[16'h041E] <= 0;
        weight_mem[16'h041F] <= 0;
        weight_mem[16'h0420] <= 0;
        weight_mem[16'h0421] <= 0;
        weight_mem[16'h0422] <= 0;
        weight_mem[16'h0423] <= 0;
        weight_mem[16'h0424] <= 0;
        weight_mem[16'h0425] <= 0;
        weight_mem[16'h0426] <= 0;
        weight_mem[16'h0427] <= 0;
        weight_mem[16'h0428] <= 0;
        weight_mem[16'h0429] <= 0;
        weight_mem[16'h042A] <= 0;
        weight_mem[16'h042B] <= 0;
        weight_mem[16'h042C] <= 0;
        weight_mem[16'h042D] <= 0;
        weight_mem[16'h042E] <= 0;
        weight_mem[16'h042F] <= 0;
        weight_mem[16'h0430] <= 0;
        weight_mem[16'h0431] <= 0;
        weight_mem[16'h0432] <= 0;
        weight_mem[16'h0433] <= 0;
        weight_mem[16'h0434] <= 0;
        weight_mem[16'h0435] <= 0;
        weight_mem[16'h0436] <= 0;
        weight_mem[16'h0437] <= 0;
        weight_mem[16'h0438] <= 0;
        weight_mem[16'h0439] <= 0;
        weight_mem[16'h043A] <= 0;
        weight_mem[16'h043B] <= 0;
        weight_mem[16'h043C] <= 0;
        weight_mem[16'h043D] <= 0;
        weight_mem[16'h043E] <= 0;
        weight_mem[16'h043F] <= 0;
        weight_mem[16'h0440] <= 0;
        weight_mem[16'h0441] <= 0;
        weight_mem[16'h0442] <= 0;
        weight_mem[16'h0443] <= 0;
        weight_mem[16'h0444] <= 0;
        weight_mem[16'h0445] <= 0;
        weight_mem[16'h0446] <= 0;
        weight_mem[16'h0447] <= 0;
        weight_mem[16'h0448] <= 0;
        weight_mem[16'h0449] <= 0;
        weight_mem[16'h044A] <= 0;
        weight_mem[16'h044B] <= 0;
        weight_mem[16'h044C] <= 0;
        weight_mem[16'h044D] <= 0;
        weight_mem[16'h044E] <= 0;
        weight_mem[16'h044F] <= 0;
        weight_mem[16'h0450] <= 0;
        weight_mem[16'h0451] <= 0;
        weight_mem[16'h0452] <= 0;
        weight_mem[16'h0453] <= 0;
        weight_mem[16'h0454] <= 0;
        weight_mem[16'h0455] <= 0;
        weight_mem[16'h0456] <= 0;
        weight_mem[16'h0457] <= 0;
        weight_mem[16'h0458] <= 0;
        weight_mem[16'h0459] <= 0;
        weight_mem[16'h045A] <= 0;
        weight_mem[16'h045B] <= 0;
        weight_mem[16'h045C] <= 0;
        weight_mem[16'h045D] <= 0;
        weight_mem[16'h045E] <= 0;
        weight_mem[16'h045F] <= 0;
        weight_mem[16'h0460] <= 0;
        weight_mem[16'h0461] <= 0;
        weight_mem[16'h0462] <= 0;
        weight_mem[16'h0463] <= 0;
        weight_mem[16'h0464] <= 0;
        weight_mem[16'h0465] <= 0;
        weight_mem[16'h0466] <= 0;
        weight_mem[16'h0467] <= 0;
        weight_mem[16'h0468] <= 0;
        weight_mem[16'h0469] <= 0;
        weight_mem[16'h046A] <= 0;
        weight_mem[16'h046B] <= 0;
        weight_mem[16'h046C] <= 0;
        weight_mem[16'h046D] <= 0;
        weight_mem[16'h046E] <= 0;
        weight_mem[16'h046F] <= 0;
        weight_mem[16'h0470] <= 0;
        weight_mem[16'h0471] <= 0;
        weight_mem[16'h0472] <= 0;
        weight_mem[16'h0473] <= 0;
        weight_mem[16'h0474] <= 0;
        weight_mem[16'h0475] <= 0;
        weight_mem[16'h0476] <= 0;
        weight_mem[16'h0477] <= 0;
        weight_mem[16'h0478] <= 0;
        weight_mem[16'h0479] <= 0;
        weight_mem[16'h047A] <= 0;
        weight_mem[16'h047B] <= 0;
        weight_mem[16'h047C] <= 0;
        weight_mem[16'h047D] <= 0;
        weight_mem[16'h047E] <= 0;
        weight_mem[16'h047F] <= 0;
        weight_mem[16'h0480] <= 0;
        weight_mem[16'h0481] <= 0;
        weight_mem[16'h0482] <= 0;
        weight_mem[16'h0483] <= 0;
        weight_mem[16'h0484] <= 0;
        weight_mem[16'h0485] <= 0;
        weight_mem[16'h0486] <= 0;
        weight_mem[16'h0487] <= 0;
        weight_mem[16'h0488] <= 0;
        weight_mem[16'h0489] <= 0;
        weight_mem[16'h048A] <= 0;
        weight_mem[16'h048B] <= 0;
        weight_mem[16'h048C] <= 0;
        weight_mem[16'h048D] <= 0;
        weight_mem[16'h048E] <= 0;
        weight_mem[16'h048F] <= 0;
        weight_mem[16'h0490] <= 0;
        weight_mem[16'h0491] <= 0;
        weight_mem[16'h0492] <= 0;
        weight_mem[16'h0493] <= 0;
        weight_mem[16'h0494] <= 0;
        weight_mem[16'h0495] <= 0;
        weight_mem[16'h0496] <= 0;
        weight_mem[16'h0497] <= 0;
        weight_mem[16'h0498] <= 0;
        weight_mem[16'h0499] <= 0;
        weight_mem[16'h049A] <= 0;
        weight_mem[16'h049B] <= 0;
        weight_mem[16'h049C] <= 0;
        weight_mem[16'h049D] <= 0;
        weight_mem[16'h049E] <= 0;
        weight_mem[16'h049F] <= 0;
        weight_mem[16'h04A0] <= 0;
        weight_mem[16'h04A1] <= 0;
        weight_mem[16'h04A2] <= 0;
        weight_mem[16'h04A3] <= 0;
        weight_mem[16'h04A4] <= 0;
        weight_mem[16'h04A5] <= 0;
        weight_mem[16'h04A6] <= 0;
        weight_mem[16'h04A7] <= 0;
        weight_mem[16'h04A8] <= 0;
        weight_mem[16'h04A9] <= 0;
        weight_mem[16'h04AA] <= 0;
        weight_mem[16'h04AB] <= 0;
        weight_mem[16'h04AC] <= 0;
        weight_mem[16'h04AD] <= 0;
        weight_mem[16'h04AE] <= 0;
        weight_mem[16'h04AF] <= 0;
        weight_mem[16'h04B0] <= 0;
        weight_mem[16'h04B1] <= 0;
        weight_mem[16'h04B2] <= 0;
        weight_mem[16'h04B3] <= 0;
        weight_mem[16'h04B4] <= 0;
        weight_mem[16'h04B5] <= 0;
        weight_mem[16'h04B6] <= 0;
        weight_mem[16'h04B7] <= 0;
        weight_mem[16'h04B8] <= 0;
        weight_mem[16'h04B9] <= 0;
        weight_mem[16'h04BA] <= 0;
        weight_mem[16'h04BB] <= 0;
        weight_mem[16'h04BC] <= 0;
        weight_mem[16'h04BD] <= 0;
        weight_mem[16'h04BE] <= 0;
        weight_mem[16'h04BF] <= 0;
        weight_mem[16'h04C0] <= 0;
        weight_mem[16'h04C1] <= 0;
        weight_mem[16'h04C2] <= 0;
        weight_mem[16'h04C3] <= 0;
        weight_mem[16'h04C4] <= 0;
        weight_mem[16'h04C5] <= 0;
        weight_mem[16'h04C6] <= 0;
        weight_mem[16'h04C7] <= 0;
        weight_mem[16'h04C8] <= 0;
        weight_mem[16'h04C9] <= 0;
        weight_mem[16'h04CA] <= 0;
        weight_mem[16'h04CB] <= 0;
        weight_mem[16'h04CC] <= 0;
        weight_mem[16'h04CD] <= 0;
        weight_mem[16'h04CE] <= 0;
        weight_mem[16'h04CF] <= 0;
        weight_mem[16'h04D0] <= 0;
        weight_mem[16'h04D1] <= 0;
        weight_mem[16'h04D2] <= 0;
        weight_mem[16'h04D3] <= 0;
        weight_mem[16'h04D4] <= 0;
        weight_mem[16'h04D5] <= 0;
        weight_mem[16'h04D6] <= 0;
        weight_mem[16'h04D7] <= 0;
        weight_mem[16'h04D8] <= 0;
        weight_mem[16'h04D9] <= 0;
        weight_mem[16'h04DA] <= 0;
        weight_mem[16'h04DB] <= 0;
        weight_mem[16'h04DC] <= 0;
        weight_mem[16'h04DD] <= 0;
        weight_mem[16'h04DE] <= 0;
        weight_mem[16'h04DF] <= 0;
        weight_mem[16'h04E0] <= 0;
        weight_mem[16'h04E1] <= 0;
        weight_mem[16'h04E2] <= 0;
        weight_mem[16'h04E3] <= 0;
        weight_mem[16'h04E4] <= 0;
        weight_mem[16'h04E5] <= 0;
        weight_mem[16'h04E6] <= 0;
        weight_mem[16'h04E7] <= 0;
        weight_mem[16'h04E8] <= 0;
        weight_mem[16'h04E9] <= 0;
        weight_mem[16'h04EA] <= 0;
        weight_mem[16'h04EB] <= 0;
        weight_mem[16'h04EC] <= 0;
        weight_mem[16'h04ED] <= 0;
        weight_mem[16'h04EE] <= 0;
        weight_mem[16'h04EF] <= 0;
        weight_mem[16'h04F0] <= 0;
        weight_mem[16'h04F1] <= 0;
        weight_mem[16'h04F2] <= 0;
        weight_mem[16'h04F3] <= 0;
        weight_mem[16'h04F4] <= 0;
        weight_mem[16'h04F5] <= 0;
        weight_mem[16'h04F6] <= 0;
        weight_mem[16'h04F7] <= 0;
        weight_mem[16'h04F8] <= 0;
        weight_mem[16'h04F9] <= 0;
        weight_mem[16'h04FA] <= 0;
        weight_mem[16'h04FB] <= 0;
        weight_mem[16'h04FC] <= 0;
        weight_mem[16'h04FD] <= 0;
        weight_mem[16'h04FE] <= 0;
        weight_mem[16'h04FF] <= 0;
        weight_mem[16'h0500] <= 0;
        weight_mem[16'h0501] <= 0;
        weight_mem[16'h0502] <= 0;
        weight_mem[16'h0503] <= 0;
        weight_mem[16'h0504] <= 0;
        weight_mem[16'h0505] <= 0;
        weight_mem[16'h0506] <= 0;
        weight_mem[16'h0507] <= 0;
        weight_mem[16'h0508] <= 0;
        weight_mem[16'h0509] <= 0;
        weight_mem[16'h050A] <= 0;
        weight_mem[16'h050B] <= 0;
        weight_mem[16'h050C] <= 0;
        weight_mem[16'h050D] <= 0;
        weight_mem[16'h050E] <= 0;
        weight_mem[16'h050F] <= 0;
        weight_mem[16'h0510] <= 0;
        weight_mem[16'h0511] <= 0;
        weight_mem[16'h0512] <= 0;
        weight_mem[16'h0513] <= 0;
        weight_mem[16'h0514] <= 0;
        weight_mem[16'h0515] <= 0;
        weight_mem[16'h0516] <= 0;
        weight_mem[16'h0517] <= 0;
        weight_mem[16'h0518] <= 0;
        weight_mem[16'h0519] <= 0;
        weight_mem[16'h051A] <= 0;
        weight_mem[16'h051B] <= 0;
        weight_mem[16'h051C] <= 0;
        weight_mem[16'h051D] <= 0;
        weight_mem[16'h051E] <= 0;
        weight_mem[16'h051F] <= 0;
        weight_mem[16'h0520] <= 0;
        weight_mem[16'h0521] <= 0;
        weight_mem[16'h0522] <= 0;
        weight_mem[16'h0523] <= 0;
        weight_mem[16'h0524] <= 0;
        weight_mem[16'h0525] <= 0;
        weight_mem[16'h0526] <= 0;
        weight_mem[16'h0527] <= 0;
        weight_mem[16'h0528] <= 0;
        weight_mem[16'h0529] <= 0;
        weight_mem[16'h052A] <= 0;
        weight_mem[16'h052B] <= 0;
        weight_mem[16'h052C] <= 0;
        weight_mem[16'h052D] <= 0;
        weight_mem[16'h052E] <= 0;
        weight_mem[16'h052F] <= 0;
        weight_mem[16'h0530] <= 0;
        weight_mem[16'h0531] <= 0;
        weight_mem[16'h0532] <= 0;
        weight_mem[16'h0533] <= 0;
        weight_mem[16'h0534] <= 0;
        weight_mem[16'h0535] <= 0;
        weight_mem[16'h0536] <= 0;
        weight_mem[16'h0537] <= 0;
        weight_mem[16'h0538] <= 0;
        weight_mem[16'h0539] <= 0;
        weight_mem[16'h053A] <= 0;
        weight_mem[16'h053B] <= 0;
        weight_mem[16'h053C] <= 0;
        weight_mem[16'h053D] <= 0;
        weight_mem[16'h053E] <= 0;
        weight_mem[16'h053F] <= 0;
        weight_mem[16'h0540] <= 0;
        weight_mem[16'h0541] <= 0;
        weight_mem[16'h0542] <= 0;
        weight_mem[16'h0543] <= 0;
        weight_mem[16'h0544] <= 0;
        weight_mem[16'h0545] <= 0;
        weight_mem[16'h0546] <= 0;
        weight_mem[16'h0547] <= 0;
        weight_mem[16'h0548] <= 0;
        weight_mem[16'h0549] <= 0;
        weight_mem[16'h054A] <= 0;
        weight_mem[16'h054B] <= 0;
        weight_mem[16'h054C] <= 0;
        weight_mem[16'h054D] <= 0;
        weight_mem[16'h054E] <= 0;
        weight_mem[16'h054F] <= 0;
        weight_mem[16'h0550] <= 0;
        weight_mem[16'h0551] <= 0;
        weight_mem[16'h0552] <= 0;
        weight_mem[16'h0553] <= 0;
        weight_mem[16'h0554] <= 0;
        weight_mem[16'h0555] <= 0;
        weight_mem[16'h0556] <= 0;
        weight_mem[16'h0557] <= 0;
        weight_mem[16'h0558] <= 0;
        weight_mem[16'h0559] <= 0;
        weight_mem[16'h055A] <= 0;
        weight_mem[16'h055B] <= 0;
        weight_mem[16'h055C] <= 0;
        weight_mem[16'h055D] <= 0;
        weight_mem[16'h055E] <= 0;
        weight_mem[16'h055F] <= 0;
        weight_mem[16'h0560] <= 0;
        weight_mem[16'h0561] <= 0;
        weight_mem[16'h0562] <= 0;
        weight_mem[16'h0563] <= 0;
        weight_mem[16'h0564] <= 0;
        weight_mem[16'h0565] <= 0;
        weight_mem[16'h0566] <= 0;
        weight_mem[16'h0567] <= 0;
        weight_mem[16'h0568] <= 0;
        weight_mem[16'h0569] <= 0;
        weight_mem[16'h056A] <= 0;
        weight_mem[16'h056B] <= 0;
        weight_mem[16'h056C] <= 0;
        weight_mem[16'h056D] <= 0;
        weight_mem[16'h056E] <= 0;
        weight_mem[16'h056F] <= 0;
        weight_mem[16'h0570] <= 0;
        weight_mem[16'h0571] <= 0;
        weight_mem[16'h0572] <= 0;
        weight_mem[16'h0573] <= 0;
        weight_mem[16'h0574] <= 0;
        weight_mem[16'h0575] <= 0;
        weight_mem[16'h0576] <= 0;
        weight_mem[16'h0577] <= 0;
        weight_mem[16'h0578] <= 0;
        weight_mem[16'h0579] <= 0;
        weight_mem[16'h057A] <= 0;
        weight_mem[16'h057B] <= 0;
        weight_mem[16'h057C] <= 0;
        weight_mem[16'h057D] <= 0;
        weight_mem[16'h057E] <= 0;
        weight_mem[16'h057F] <= 0;
        weight_mem[16'h0580] <= 0;
        weight_mem[16'h0581] <= 0;
        weight_mem[16'h0582] <= 0;
        weight_mem[16'h0583] <= 0;
        weight_mem[16'h0584] <= 0;
        weight_mem[16'h0585] <= 0;
        weight_mem[16'h0586] <= 0;
        weight_mem[16'h0587] <= 0;
        weight_mem[16'h0588] <= 0;
        weight_mem[16'h0589] <= 0;
        weight_mem[16'h058A] <= 0;
        weight_mem[16'h058B] <= 0;
        weight_mem[16'h058C] <= 0;
        weight_mem[16'h058D] <= 0;
        weight_mem[16'h058E] <= 0;
        weight_mem[16'h058F] <= 0;
        weight_mem[16'h0590] <= 0;
        weight_mem[16'h0591] <= 0;
        weight_mem[16'h0592] <= 0;
        weight_mem[16'h0593] <= 0;
        weight_mem[16'h0594] <= 0;
        weight_mem[16'h0595] <= 0;
        weight_mem[16'h0596] <= 0;
        weight_mem[16'h0597] <= 0;
        weight_mem[16'h0598] <= 0;
        weight_mem[16'h0599] <= 0;
        weight_mem[16'h059A] <= 0;
        weight_mem[16'h059B] <= 0;
        weight_mem[16'h059C] <= 0;
        weight_mem[16'h059D] <= 0;
        weight_mem[16'h059E] <= 0;
        weight_mem[16'h059F] <= 0;
        weight_mem[16'h05A0] <= 0;
        weight_mem[16'h05A1] <= 0;
        weight_mem[16'h05A2] <= 0;
        weight_mem[16'h05A3] <= 0;
        weight_mem[16'h05A4] <= 0;
        weight_mem[16'h05A5] <= 0;
        weight_mem[16'h05A6] <= 0;
        weight_mem[16'h05A7] <= 0;
        weight_mem[16'h05A8] <= 0;
        weight_mem[16'h05A9] <= 0;
        weight_mem[16'h05AA] <= 0;
        weight_mem[16'h05AB] <= 0;
        weight_mem[16'h05AC] <= 0;
        weight_mem[16'h05AD] <= 0;
        weight_mem[16'h05AE] <= 0;
        weight_mem[16'h05AF] <= 0;

        // layer 1 neuron 3
        weight_mem[16'h0600] <= 0;
        weight_mem[16'h0601] <= 0;
        weight_mem[16'h0602] <= 0;
        weight_mem[16'h0603] <= 0;
        weight_mem[16'h0604] <= 0;
        weight_mem[16'h0605] <= 0;
        weight_mem[16'h0606] <= 0;
        weight_mem[16'h0607] <= 0;
        weight_mem[16'h0608] <= 0;
        weight_mem[16'h0609] <= 0;
        weight_mem[16'h060A] <= 0;
        weight_mem[16'h060B] <= 0;
        weight_mem[16'h060C] <= 0;
        weight_mem[16'h060D] <= 0;
        weight_mem[16'h060E] <= 0;
        weight_mem[16'h060F] <= 0;
        weight_mem[16'h0610] <= 0;
        weight_mem[16'h0611] <= 0;
        weight_mem[16'h0612] <= 0;
        weight_mem[16'h0613] <= 0;
        weight_mem[16'h0614] <= 0;
        weight_mem[16'h0615] <= 0;
        weight_mem[16'h0616] <= 0;
        weight_mem[16'h0617] <= 0;
        weight_mem[16'h0618] <= 0;
        weight_mem[16'h0619] <= 0;
        weight_mem[16'h061A] <= 0;
        weight_mem[16'h061B] <= 0;
        weight_mem[16'h061C] <= 0;
        weight_mem[16'h061D] <= 0;
        weight_mem[16'h061E] <= 0;
        weight_mem[16'h061F] <= 0;
        weight_mem[16'h0620] <= 0;
        weight_mem[16'h0621] <= 0;
        weight_mem[16'h0622] <= 0;
        weight_mem[16'h0623] <= 0;
        weight_mem[16'h0624] <= 0;
        weight_mem[16'h0625] <= 0;
        weight_mem[16'h0626] <= 0;
        weight_mem[16'h0627] <= 0;
        weight_mem[16'h0628] <= 0;
        weight_mem[16'h0629] <= 0;
        weight_mem[16'h062A] <= 0;
        weight_mem[16'h062B] <= 0;
        weight_mem[16'h062C] <= 0;
        weight_mem[16'h062D] <= 0;
        weight_mem[16'h062E] <= 0;
        weight_mem[16'h062F] <= 0;
        weight_mem[16'h0630] <= 0;
        weight_mem[16'h0631] <= 0;
        weight_mem[16'h0632] <= 0;
        weight_mem[16'h0633] <= 0;
        weight_mem[16'h0634] <= 0;
        weight_mem[16'h0635] <= 0;
        weight_mem[16'h0636] <= 0;
        weight_mem[16'h0637] <= 0;
        weight_mem[16'h0638] <= 0;
        weight_mem[16'h0639] <= 0;
        weight_mem[16'h063A] <= 0;
        weight_mem[16'h063B] <= 0;
        weight_mem[16'h063C] <= 0;
        weight_mem[16'h063D] <= 0;
        weight_mem[16'h063E] <= 0;
        weight_mem[16'h063F] <= 0;
        weight_mem[16'h0640] <= 0;
        weight_mem[16'h0641] <= 0;
        weight_mem[16'h0642] <= 0;
        weight_mem[16'h0643] <= 0;
        weight_mem[16'h0644] <= 0;
        weight_mem[16'h0645] <= 0;
        weight_mem[16'h0646] <= 0;
        weight_mem[16'h0647] <= 0;
        weight_mem[16'h0648] <= 0;
        weight_mem[16'h0649] <= 0;
        weight_mem[16'h064A] <= 0;
        weight_mem[16'h064B] <= 0;
        weight_mem[16'h064C] <= 0;
        weight_mem[16'h064D] <= 0;
        weight_mem[16'h064E] <= 0;
        weight_mem[16'h064F] <= 0;
        weight_mem[16'h0650] <= 0;
        weight_mem[16'h0651] <= 0;
        weight_mem[16'h0652] <= 0;
        weight_mem[16'h0653] <= 0;
        weight_mem[16'h0654] <= 0;
        weight_mem[16'h0655] <= 0;
        weight_mem[16'h0656] <= 0;
        weight_mem[16'h0657] <= 0;
        weight_mem[16'h0658] <= 0;
        weight_mem[16'h0659] <= 0;
        weight_mem[16'h065A] <= 0;
        weight_mem[16'h065B] <= 0;
        weight_mem[16'h065C] <= 0;
        weight_mem[16'h065D] <= 0;
        weight_mem[16'h065E] <= 0;
        weight_mem[16'h065F] <= 0;
        weight_mem[16'h0660] <= 0;
        weight_mem[16'h0661] <= 0;
        weight_mem[16'h0662] <= 0;
        weight_mem[16'h0663] <= 0;
        weight_mem[16'h0664] <= 0;
        weight_mem[16'h0665] <= 0;
        weight_mem[16'h0666] <= 0;
        weight_mem[16'h0667] <= 0;
        weight_mem[16'h0668] <= 0;
        weight_mem[16'h0669] <= 0;
        weight_mem[16'h066A] <= 0;
        weight_mem[16'h066B] <= 0;
        weight_mem[16'h066C] <= 0;
        weight_mem[16'h066D] <= 0;
        weight_mem[16'h066E] <= 0;
        weight_mem[16'h066F] <= 0;
        weight_mem[16'h0670] <= 0;
        weight_mem[16'h0671] <= 0;
        weight_mem[16'h0672] <= 0;
        weight_mem[16'h0673] <= 0;
        weight_mem[16'h0674] <= 0;
        weight_mem[16'h0675] <= 0;
        weight_mem[16'h0676] <= 0;
        weight_mem[16'h0677] <= 0;
        weight_mem[16'h0678] <= 0;
        weight_mem[16'h0679] <= 0;
        weight_mem[16'h067A] <= 0;
        weight_mem[16'h067B] <= 0;
        weight_mem[16'h067C] <= 0;
        weight_mem[16'h067D] <= 0;
        weight_mem[16'h067E] <= 0;
        weight_mem[16'h067F] <= 0;
        weight_mem[16'h0680] <= 0;
        weight_mem[16'h0681] <= 0;
        weight_mem[16'h0682] <= 0;
        weight_mem[16'h0683] <= 0;
        weight_mem[16'h0684] <= 0;
        weight_mem[16'h0685] <= 0;
        weight_mem[16'h0686] <= 0;
        weight_mem[16'h0687] <= 0;
        weight_mem[16'h0688] <= 0;
        weight_mem[16'h0689] <= 0;
        weight_mem[16'h068A] <= 0;
        weight_mem[16'h068B] <= 0;
        weight_mem[16'h068C] <= 0;
        weight_mem[16'h068D] <= 0;
        weight_mem[16'h068E] <= 0;
        weight_mem[16'h068F] <= 0;
        weight_mem[16'h0690] <= 0;
        weight_mem[16'h0691] <= 0;
        weight_mem[16'h0692] <= 0;
        weight_mem[16'h0693] <= 0;
        weight_mem[16'h0694] <= 0;
        weight_mem[16'h0695] <= 0;
        weight_mem[16'h0696] <= 0;
        weight_mem[16'h0697] <= 0;
        weight_mem[16'h0698] <= 0;
        weight_mem[16'h0699] <= 0;
        weight_mem[16'h069A] <= 0;
        weight_mem[16'h069B] <= 0;
        weight_mem[16'h069C] <= 0;
        weight_mem[16'h069D] <= 0;
        weight_mem[16'h069E] <= 0;
        weight_mem[16'h069F] <= 0;
        weight_mem[16'h06A0] <= 0;
        weight_mem[16'h06A1] <= 0;
        weight_mem[16'h06A2] <= 0;
        weight_mem[16'h06A3] <= 0;
        weight_mem[16'h06A4] <= 0;
        weight_mem[16'h06A5] <= 0;
        weight_mem[16'h06A6] <= 0;
        weight_mem[16'h06A7] <= 0;
        weight_mem[16'h06A8] <= 0;
        weight_mem[16'h06A9] <= 0;
        weight_mem[16'h06AA] <= 0;
        weight_mem[16'h06AB] <= 0;
        weight_mem[16'h06AC] <= 0;
        weight_mem[16'h06AD] <= 0;
        weight_mem[16'h06AE] <= 0;
        weight_mem[16'h06AF] <= 0;
        weight_mem[16'h06B0] <= 0;
        weight_mem[16'h06B1] <= 0;
        weight_mem[16'h06B2] <= 0;
        weight_mem[16'h06B3] <= 0;
        weight_mem[16'h06B4] <= 0;
        weight_mem[16'h06B5] <= 0;
        weight_mem[16'h06B6] <= 0;
        weight_mem[16'h06B7] <= 0;
        weight_mem[16'h06B8] <= 0;
        weight_mem[16'h06B9] <= 0;
        weight_mem[16'h06BA] <= 0;
        weight_mem[16'h06BB] <= 0;
        weight_mem[16'h06BC] <= 0;
        weight_mem[16'h06BD] <= 0;
        weight_mem[16'h06BE] <= 0;
        weight_mem[16'h06BF] <= 0;
        weight_mem[16'h06C0] <= 0;
        weight_mem[16'h06C1] <= 0;
        weight_mem[16'h06C2] <= 0;
        weight_mem[16'h06C3] <= 0;
        weight_mem[16'h06C4] <= 0;
        weight_mem[16'h06C5] <= 0;
        weight_mem[16'h06C6] <= 0;
        weight_mem[16'h06C7] <= 0;
        weight_mem[16'h06C8] <= 0;
        weight_mem[16'h06C9] <= 0;
        weight_mem[16'h06CA] <= 0;
        weight_mem[16'h06CB] <= 0;
        weight_mem[16'h06CC] <= 0;
        weight_mem[16'h06CD] <= 0;
        weight_mem[16'h06CE] <= 0;
        weight_mem[16'h06CF] <= 0;
        weight_mem[16'h06D0] <= 0;
        weight_mem[16'h06D1] <= 0;
        weight_mem[16'h06D2] <= 0;
        weight_mem[16'h06D3] <= 0;
        weight_mem[16'h06D4] <= 0;
        weight_mem[16'h06D5] <= 0;
        weight_mem[16'h06D6] <= 0;
        weight_mem[16'h06D7] <= 0;
        weight_mem[16'h06D8] <= 0;
        weight_mem[16'h06D9] <= 0;
        weight_mem[16'h06DA] <= 0;
        weight_mem[16'h06DB] <= 0;
        weight_mem[16'h06DC] <= 0;
        weight_mem[16'h06DD] <= 0;
        weight_mem[16'h06DE] <= 0;
        weight_mem[16'h06DF] <= 0;
        weight_mem[16'h06E0] <= 0;
        weight_mem[16'h06E1] <= 0;
        weight_mem[16'h06E2] <= 0;
        weight_mem[16'h06E3] <= 0;
        weight_mem[16'h06E4] <= 0;
        weight_mem[16'h06E5] <= 0;
        weight_mem[16'h06E6] <= 0;
        weight_mem[16'h06E7] <= 0;
        weight_mem[16'h06E8] <= 0;
        weight_mem[16'h06E9] <= 0;
        weight_mem[16'h06EA] <= 0;
        weight_mem[16'h06EB] <= 0;
        weight_mem[16'h06EC] <= 0;
        weight_mem[16'h06ED] <= 0;
        weight_mem[16'h06EE] <= 0;
        weight_mem[16'h06EF] <= 0;
        weight_mem[16'h06F0] <= 0;
        weight_mem[16'h06F1] <= 0;
        weight_mem[16'h06F2] <= 0;
        weight_mem[16'h06F3] <= 0;
        weight_mem[16'h06F4] <= 0;
        weight_mem[16'h06F5] <= 0;
        weight_mem[16'h06F6] <= 0;
        weight_mem[16'h06F7] <= 0;
        weight_mem[16'h06F8] <= 0;
        weight_mem[16'h06F9] <= 0;
        weight_mem[16'h06FA] <= 0;
        weight_mem[16'h06FB] <= 0;
        weight_mem[16'h06FC] <= 0;
        weight_mem[16'h06FD] <= 0;
        weight_mem[16'h06FE] <= 0;
        weight_mem[16'h06FF] <= 0;
        weight_mem[16'h0700] <= 0;
        weight_mem[16'h0701] <= 0;
        weight_mem[16'h0702] <= 0;
        weight_mem[16'h0703] <= 0;
        weight_mem[16'h0704] <= 0;
        weight_mem[16'h0705] <= 0;
        weight_mem[16'h0706] <= 0;
        weight_mem[16'h0707] <= 0;
        weight_mem[16'h0708] <= 0;
        weight_mem[16'h0709] <= 0;
        weight_mem[16'h070A] <= 0;
        weight_mem[16'h070B] <= 0;
        weight_mem[16'h070C] <= 0;
        weight_mem[16'h070D] <= 0;
        weight_mem[16'h070E] <= 0;
        weight_mem[16'h070F] <= 0;
        weight_mem[16'h0710] <= 0;
        weight_mem[16'h0711] <= 0;
        weight_mem[16'h0712] <= 0;
        weight_mem[16'h0713] <= 0;
        weight_mem[16'h0714] <= 0;
        weight_mem[16'h0715] <= 0;
        weight_mem[16'h0716] <= 0;
        weight_mem[16'h0717] <= 0;
        weight_mem[16'h0718] <= 0;
        weight_mem[16'h0719] <= 0;
        weight_mem[16'h071A] <= 0;
        weight_mem[16'h071B] <= 0;
        weight_mem[16'h071C] <= 0;
        weight_mem[16'h071D] <= 0;
        weight_mem[16'h071E] <= 0;
        weight_mem[16'h071F] <= 0;
        weight_mem[16'h0720] <= 0;
        weight_mem[16'h0721] <= 0;
        weight_mem[16'h0722] <= 0;
        weight_mem[16'h0723] <= 0;
        weight_mem[16'h0724] <= 0;
        weight_mem[16'h0725] <= 0;
        weight_mem[16'h0726] <= 0;
        weight_mem[16'h0727] <= 0;
        weight_mem[16'h0728] <= 0;
        weight_mem[16'h0729] <= 0;
        weight_mem[16'h072A] <= 0;
        weight_mem[16'h072B] <= 0;
        weight_mem[16'h072C] <= 0;
        weight_mem[16'h072D] <= 0;
        weight_mem[16'h072E] <= 0;
        weight_mem[16'h072F] <= 0;
        weight_mem[16'h0730] <= 0;
        weight_mem[16'h0731] <= 0;
        weight_mem[16'h0732] <= 0;
        weight_mem[16'h0733] <= 0;
        weight_mem[16'h0734] <= 0;
        weight_mem[16'h0735] <= 0;
        weight_mem[16'h0736] <= 0;
        weight_mem[16'h0737] <= 0;
        weight_mem[16'h0738] <= 0;
        weight_mem[16'h0739] <= 0;
        weight_mem[16'h073A] <= 0;
        weight_mem[16'h073B] <= 0;
        weight_mem[16'h073C] <= 0;
        weight_mem[16'h073D] <= 0;
        weight_mem[16'h073E] <= 0;
        weight_mem[16'h073F] <= 0;
        weight_mem[16'h0740] <= 0;
        weight_mem[16'h0741] <= 0;
        weight_mem[16'h0742] <= 0;
        weight_mem[16'h0743] <= 0;
        weight_mem[16'h0744] <= 0;
        weight_mem[16'h0745] <= 0;
        weight_mem[16'h0746] <= 0;
        weight_mem[16'h0747] <= 0;
        weight_mem[16'h0748] <= 0;
        weight_mem[16'h0749] <= 0;
        weight_mem[16'h074A] <= 0;
        weight_mem[16'h074B] <= 0;
        weight_mem[16'h074C] <= 0;
        weight_mem[16'h074D] <= 0;
        weight_mem[16'h074E] <= 0;
        weight_mem[16'h074F] <= 0;
        weight_mem[16'h0750] <= 0;
        weight_mem[16'h0751] <= 0;
        weight_mem[16'h0752] <= 0;
        weight_mem[16'h0753] <= 0;
        weight_mem[16'h0754] <= 0;
        weight_mem[16'h0755] <= 0;
        weight_mem[16'h0756] <= 0;
        weight_mem[16'h0757] <= 0;
        weight_mem[16'h0758] <= 0;
        weight_mem[16'h0759] <= 0;
        weight_mem[16'h075A] <= 0;
        weight_mem[16'h075B] <= 0;
        weight_mem[16'h075C] <= 0;
        weight_mem[16'h075D] <= 0;
        weight_mem[16'h075E] <= 0;
        weight_mem[16'h075F] <= 0;
        weight_mem[16'h0760] <= 0;
        weight_mem[16'h0761] <= 0;
        weight_mem[16'h0762] <= 0;
        weight_mem[16'h0763] <= 0;
        weight_mem[16'h0764] <= 0;
        weight_mem[16'h0765] <= 0;
        weight_mem[16'h0766] <= 0;
        weight_mem[16'h0767] <= 0;
        weight_mem[16'h0768] <= 0;
        weight_mem[16'h0769] <= 0;
        weight_mem[16'h076A] <= 0;
        weight_mem[16'h076B] <= 0;
        weight_mem[16'h076C] <= 0;
        weight_mem[16'h076D] <= 0;
        weight_mem[16'h076E] <= 0;
        weight_mem[16'h076F] <= 0;
        weight_mem[16'h0770] <= 0;
        weight_mem[16'h0771] <= 0;
        weight_mem[16'h0772] <= 0;
        weight_mem[16'h0773] <= 0;
        weight_mem[16'h0774] <= 0;
        weight_mem[16'h0775] <= 0;
        weight_mem[16'h0776] <= 0;
        weight_mem[16'h0777] <= 0;
        weight_mem[16'h0778] <= 0;
        weight_mem[16'h0779] <= 0;
        weight_mem[16'h077A] <= 0;
        weight_mem[16'h077B] <= 0;
        weight_mem[16'h077C] <= 0;
        weight_mem[16'h077D] <= 0;
        weight_mem[16'h077E] <= 0;
        weight_mem[16'h077F] <= 0;
        weight_mem[16'h0780] <= 0;
        weight_mem[16'h0781] <= 0;
        weight_mem[16'h0782] <= 0;
        weight_mem[16'h0783] <= 0;
        weight_mem[16'h0784] <= 0;
        weight_mem[16'h0785] <= 0;
        weight_mem[16'h0786] <= 0;
        weight_mem[16'h0787] <= 0;
        weight_mem[16'h0788] <= 0;
        weight_mem[16'h0789] <= 0;
        weight_mem[16'h078A] <= 0;
        weight_mem[16'h078B] <= 0;
        weight_mem[16'h078C] <= 0;
        weight_mem[16'h078D] <= 0;
        weight_mem[16'h078E] <= 0;
        weight_mem[16'h078F] <= 0;
        weight_mem[16'h0790] <= 0;
        weight_mem[16'h0791] <= 0;
        weight_mem[16'h0792] <= 0;
        weight_mem[16'h0793] <= 0;
        weight_mem[16'h0794] <= 0;
        weight_mem[16'h0795] <= 0;
        weight_mem[16'h0796] <= 0;
        weight_mem[16'h0797] <= 0;
        weight_mem[16'h0798] <= 0;
        weight_mem[16'h0799] <= 0;
        weight_mem[16'h079A] <= 0;
        weight_mem[16'h079B] <= 0;
        weight_mem[16'h079C] <= 0;
        weight_mem[16'h079D] <= 0;
        weight_mem[16'h079E] <= 0;
        weight_mem[16'h079F] <= 0;
        weight_mem[16'h07A0] <= 0;
        weight_mem[16'h07A1] <= 0;
        weight_mem[16'h07A2] <= 0;
        weight_mem[16'h07A3] <= 0;
        weight_mem[16'h07A4] <= 0;
        weight_mem[16'h07A5] <= 0;
        weight_mem[16'h07A6] <= 0;
        weight_mem[16'h07A7] <= 0;
        weight_mem[16'h07A8] <= 0;
        weight_mem[16'h07A9] <= 0;
        weight_mem[16'h07AA] <= 0;
        weight_mem[16'h07AB] <= 0;
        weight_mem[16'h07AC] <= 0;
        weight_mem[16'h07AD] <= 0;
        weight_mem[16'h07AE] <= 0;
        weight_mem[16'h07AF] <= 0;

        // layer 1 neuron 4
        weight_mem[16'h0800] <= 0;
        weight_mem[16'h0801] <= 0;
        weight_mem[16'h0802] <= 0;
        weight_mem[16'h0803] <= 0;
        weight_mem[16'h0804] <= 0;
        weight_mem[16'h0805] <= 0;
        weight_mem[16'h0806] <= 0;
        weight_mem[16'h0807] <= 0;
        weight_mem[16'h0808] <= 0;
        weight_mem[16'h0809] <= 0;
        weight_mem[16'h080A] <= 0;
        weight_mem[16'h080B] <= 0;
        weight_mem[16'h080C] <= 0;
        weight_mem[16'h080D] <= 0;
        weight_mem[16'h080E] <= 0;
        weight_mem[16'h080F] <= 0;
        weight_mem[16'h0810] <= 0;
        weight_mem[16'h0811] <= 0;
        weight_mem[16'h0812] <= 0;
        weight_mem[16'h0813] <= 0;
        weight_mem[16'h0814] <= 0;
        weight_mem[16'h0815] <= 0;
        weight_mem[16'h0816] <= 0;
        weight_mem[16'h0817] <= 0;
        weight_mem[16'h0818] <= 0;
        weight_mem[16'h0819] <= 0;
        weight_mem[16'h081A] <= 0;
        weight_mem[16'h081B] <= 0;
        weight_mem[16'h081C] <= 0;
        weight_mem[16'h081D] <= 0;
        weight_mem[16'h081E] <= 0;
        weight_mem[16'h081F] <= 0;
        weight_mem[16'h0820] <= 0;
        weight_mem[16'h0821] <= 0;
        weight_mem[16'h0822] <= 0;
        weight_mem[16'h0823] <= 0;
        weight_mem[16'h0824] <= 0;
        weight_mem[16'h0825] <= 0;
        weight_mem[16'h0826] <= 0;
        weight_mem[16'h0827] <= 0;
        weight_mem[16'h0828] <= 0;
        weight_mem[16'h0829] <= 0;
        weight_mem[16'h082A] <= 0;
        weight_mem[16'h082B] <= 0;
        weight_mem[16'h082C] <= 0;
        weight_mem[16'h082D] <= 0;
        weight_mem[16'h082E] <= 0;
        weight_mem[16'h082F] <= 0;
        weight_mem[16'h0830] <= 0;
        weight_mem[16'h0831] <= 0;
        weight_mem[16'h0832] <= 0;
        weight_mem[16'h0833] <= 0;
        weight_mem[16'h0834] <= 0;
        weight_mem[16'h0835] <= 0;
        weight_mem[16'h0836] <= 0;
        weight_mem[16'h0837] <= 0;
        weight_mem[16'h0838] <= 0;
        weight_mem[16'h0839] <= 0;
        weight_mem[16'h083A] <= 0;
        weight_mem[16'h083B] <= 0;
        weight_mem[16'h083C] <= 0;
        weight_mem[16'h083D] <= 0;
        weight_mem[16'h083E] <= 0;
        weight_mem[16'h083F] <= 0;
        weight_mem[16'h0840] <= 0;
        weight_mem[16'h0841] <= 0;
        weight_mem[16'h0842] <= 0;
        weight_mem[16'h0843] <= 0;
        weight_mem[16'h0844] <= 0;
        weight_mem[16'h0845] <= 0;
        weight_mem[16'h0846] <= 0;
        weight_mem[16'h0847] <= 0;
        weight_mem[16'h0848] <= 0;
        weight_mem[16'h0849] <= 0;
        weight_mem[16'h084A] <= 0;
        weight_mem[16'h084B] <= 0;
        weight_mem[16'h084C] <= 0;
        weight_mem[16'h084D] <= 0;
        weight_mem[16'h084E] <= 0;
        weight_mem[16'h084F] <= 0;
        weight_mem[16'h0850] <= 0;
        weight_mem[16'h0851] <= 0;
        weight_mem[16'h0852] <= 0;
        weight_mem[16'h0853] <= 0;
        weight_mem[16'h0854] <= 0;
        weight_mem[16'h0855] <= 0;
        weight_mem[16'h0856] <= 0;
        weight_mem[16'h0857] <= 0;
        weight_mem[16'h0858] <= 0;
        weight_mem[16'h0859] <= 0;
        weight_mem[16'h085A] <= 0;
        weight_mem[16'h085B] <= 0;
        weight_mem[16'h085C] <= 0;
        weight_mem[16'h085D] <= 0;
        weight_mem[16'h085E] <= 0;
        weight_mem[16'h085F] <= 0;
        weight_mem[16'h0860] <= 0;
        weight_mem[16'h0861] <= 0;
        weight_mem[16'h0862] <= 0;
        weight_mem[16'h0863] <= 0;
        weight_mem[16'h0864] <= 0;
        weight_mem[16'h0865] <= 0;
        weight_mem[16'h0866] <= 0;
        weight_mem[16'h0867] <= 0;
        weight_mem[16'h0868] <= 0;
        weight_mem[16'h0869] <= 0;
        weight_mem[16'h086A] <= 0;
        weight_mem[16'h086B] <= 0;
        weight_mem[16'h086C] <= 0;
        weight_mem[16'h086D] <= 0;
        weight_mem[16'h086E] <= 0;
        weight_mem[16'h086F] <= 0;
        weight_mem[16'h0870] <= 0;
        weight_mem[16'h0871] <= 0;
        weight_mem[16'h0872] <= 0;
        weight_mem[16'h0873] <= 0;
        weight_mem[16'h0874] <= 0;
        weight_mem[16'h0875] <= 0;
        weight_mem[16'h0876] <= 0;
        weight_mem[16'h0877] <= 0;
        weight_mem[16'h0878] <= 0;
        weight_mem[16'h0879] <= 0;
        weight_mem[16'h087A] <= 0;
        weight_mem[16'h087B] <= 0;
        weight_mem[16'h087C] <= 0;
        weight_mem[16'h087D] <= 0;
        weight_mem[16'h087E] <= 0;
        weight_mem[16'h087F] <= 0;
        weight_mem[16'h0880] <= 0;
        weight_mem[16'h0881] <= 0;
        weight_mem[16'h0882] <= 0;
        weight_mem[16'h0883] <= 0;
        weight_mem[16'h0884] <= 0;
        weight_mem[16'h0885] <= 0;
        weight_mem[16'h0886] <= 0;
        weight_mem[16'h0887] <= 0;
        weight_mem[16'h0888] <= 0;
        weight_mem[16'h0889] <= 0;
        weight_mem[16'h088A] <= 0;
        weight_mem[16'h088B] <= 0;
        weight_mem[16'h088C] <= 0;
        weight_mem[16'h088D] <= 0;
        weight_mem[16'h088E] <= 0;
        weight_mem[16'h088F] <= 0;
        weight_mem[16'h0890] <= 0;
        weight_mem[16'h0891] <= 0;
        weight_mem[16'h0892] <= 0;
        weight_mem[16'h0893] <= 0;
        weight_mem[16'h0894] <= 0;
        weight_mem[16'h0895] <= 0;
        weight_mem[16'h0896] <= 0;
        weight_mem[16'h0897] <= 0;
        weight_mem[16'h0898] <= 0;
        weight_mem[16'h0899] <= 0;
        weight_mem[16'h089A] <= 0;
        weight_mem[16'h089B] <= 0;
        weight_mem[16'h089C] <= 0;
        weight_mem[16'h089D] <= 0;
        weight_mem[16'h089E] <= 0;
        weight_mem[16'h089F] <= 0;
        weight_mem[16'h08A0] <= 0;
        weight_mem[16'h08A1] <= 0;
        weight_mem[16'h08A2] <= 0;
        weight_mem[16'h08A3] <= 0;
        weight_mem[16'h08A4] <= 0;
        weight_mem[16'h08A5] <= 0;
        weight_mem[16'h08A6] <= 0;
        weight_mem[16'h08A7] <= 0;
        weight_mem[16'h08A8] <= 0;
        weight_mem[16'h08A9] <= 0;
        weight_mem[16'h08AA] <= 0;
        weight_mem[16'h08AB] <= 0;
        weight_mem[16'h08AC] <= 0;
        weight_mem[16'h08AD] <= 0;
        weight_mem[16'h08AE] <= 0;
        weight_mem[16'h08AF] <= 0;
        weight_mem[16'h08B0] <= 0;
        weight_mem[16'h08B1] <= 0;
        weight_mem[16'h08B2] <= 0;
        weight_mem[16'h08B3] <= 0;
        weight_mem[16'h08B4] <= 0;
        weight_mem[16'h08B5] <= 0;
        weight_mem[16'h08B6] <= 0;
        weight_mem[16'h08B7] <= 0;
        weight_mem[16'h08B8] <= 0;
        weight_mem[16'h08B9] <= 0;
        weight_mem[16'h08BA] <= 0;
        weight_mem[16'h08BB] <= 0;
        weight_mem[16'h08BC] <= 0;
        weight_mem[16'h08BD] <= 0;
        weight_mem[16'h08BE] <= 0;
        weight_mem[16'h08BF] <= 0;
        weight_mem[16'h08C0] <= 0;
        weight_mem[16'h08C1] <= 0;
        weight_mem[16'h08C2] <= 0;
        weight_mem[16'h08C3] <= 0;
        weight_mem[16'h08C4] <= 0;
        weight_mem[16'h08C5] <= 0;
        weight_mem[16'h08C6] <= 0;
        weight_mem[16'h08C7] <= 0;
        weight_mem[16'h08C8] <= 0;
        weight_mem[16'h08C9] <= 0;
        weight_mem[16'h08CA] <= 0;
        weight_mem[16'h08CB] <= 0;
        weight_mem[16'h08CC] <= 0;
        weight_mem[16'h08CD] <= 0;
        weight_mem[16'h08CE] <= 0;
        weight_mem[16'h08CF] <= 0;
        weight_mem[16'h08D0] <= 0;
        weight_mem[16'h08D1] <= 0;
        weight_mem[16'h08D2] <= 0;
        weight_mem[16'h08D3] <= 0;
        weight_mem[16'h08D4] <= 0;
        weight_mem[16'h08D5] <= 0;
        weight_mem[16'h08D6] <= 0;
        weight_mem[16'h08D7] <= 0;
        weight_mem[16'h08D8] <= 0;
        weight_mem[16'h08D9] <= 0;
        weight_mem[16'h08DA] <= 0;
        weight_mem[16'h08DB] <= 0;
        weight_mem[16'h08DC] <= 0;
        weight_mem[16'h08DD] <= 0;
        weight_mem[16'h08DE] <= 0;
        weight_mem[16'h08DF] <= 0;
        weight_mem[16'h08E0] <= 0;
        weight_mem[16'h08E1] <= 0;
        weight_mem[16'h08E2] <= 0;
        weight_mem[16'h08E3] <= 0;
        weight_mem[16'h08E4] <= 0;
        weight_mem[16'h08E5] <= 0;
        weight_mem[16'h08E6] <= 0;
        weight_mem[16'h08E7] <= 0;
        weight_mem[16'h08E8] <= 0;
        weight_mem[16'h08E9] <= 0;
        weight_mem[16'h08EA] <= 0;
        weight_mem[16'h08EB] <= 0;
        weight_mem[16'h08EC] <= 0;
        weight_mem[16'h08ED] <= 0;
        weight_mem[16'h08EE] <= 0;
        weight_mem[16'h08EF] <= 0;
        weight_mem[16'h08F0] <= 0;
        weight_mem[16'h08F1] <= 0;
        weight_mem[16'h08F2] <= 0;
        weight_mem[16'h08F3] <= 0;
        weight_mem[16'h08F4] <= 0;
        weight_mem[16'h08F5] <= 0;
        weight_mem[16'h08F6] <= 0;
        weight_mem[16'h08F7] <= 0;
        weight_mem[16'h08F8] <= 0;
        weight_mem[16'h08F9] <= 0;
        weight_mem[16'h08FA] <= 0;
        weight_mem[16'h08FB] <= 0;
        weight_mem[16'h08FC] <= 0;
        weight_mem[16'h08FD] <= 0;
        weight_mem[16'h08FE] <= 0;
        weight_mem[16'h08FF] <= 0;
        weight_mem[16'h0900] <= 0;
        weight_mem[16'h0901] <= 0;
        weight_mem[16'h0902] <= 0;
        weight_mem[16'h0903] <= 0;
        weight_mem[16'h0904] <= 0;
        weight_mem[16'h0905] <= 0;
        weight_mem[16'h0906] <= 0;
        weight_mem[16'h0907] <= 0;
        weight_mem[16'h0908] <= 0;
        weight_mem[16'h0909] <= 0;
        weight_mem[16'h090A] <= 0;
        weight_mem[16'h090B] <= 0;
        weight_mem[16'h090C] <= 0;
        weight_mem[16'h090D] <= 0;
        weight_mem[16'h090E] <= 0;
        weight_mem[16'h090F] <= 0;
        weight_mem[16'h0910] <= 0;
        weight_mem[16'h0911] <= 0;
        weight_mem[16'h0912] <= 0;
        weight_mem[16'h0913] <= 0;
        weight_mem[16'h0914] <= 0;
        weight_mem[16'h0915] <= 0;
        weight_mem[16'h0916] <= 0;
        weight_mem[16'h0917] <= 0;
        weight_mem[16'h0918] <= 0;
        weight_mem[16'h0919] <= 0;
        weight_mem[16'h091A] <= 0;
        weight_mem[16'h091B] <= 0;
        weight_mem[16'h091C] <= 0;
        weight_mem[16'h091D] <= 0;
        weight_mem[16'h091E] <= 0;
        weight_mem[16'h091F] <= 0;
        weight_mem[16'h0920] <= 0;
        weight_mem[16'h0921] <= 0;
        weight_mem[16'h0922] <= 0;
        weight_mem[16'h0923] <= 0;
        weight_mem[16'h0924] <= 0;
        weight_mem[16'h0925] <= 0;
        weight_mem[16'h0926] <= 0;
        weight_mem[16'h0927] <= 0;
        weight_mem[16'h0928] <= 0;
        weight_mem[16'h0929] <= 0;
        weight_mem[16'h092A] <= 0;
        weight_mem[16'h092B] <= 0;
        weight_mem[16'h092C] <= 0;
        weight_mem[16'h092D] <= 0;
        weight_mem[16'h092E] <= 0;
        weight_mem[16'h092F] <= 0;
        weight_mem[16'h0930] <= 0;
        weight_mem[16'h0931] <= 0;
        weight_mem[16'h0932] <= 0;
        weight_mem[16'h0933] <= 0;
        weight_mem[16'h0934] <= 0;
        weight_mem[16'h0935] <= 0;
        weight_mem[16'h0936] <= 0;
        weight_mem[16'h0937] <= 0;
        weight_mem[16'h0938] <= 0;
        weight_mem[16'h0939] <= 0;
        weight_mem[16'h093A] <= 0;
        weight_mem[16'h093B] <= 0;
        weight_mem[16'h093C] <= 0;
        weight_mem[16'h093D] <= 0;
        weight_mem[16'h093E] <= 0;
        weight_mem[16'h093F] <= 0;
        weight_mem[16'h0940] <= 0;
        weight_mem[16'h0941] <= 0;
        weight_mem[16'h0942] <= 0;
        weight_mem[16'h0943] <= 0;
        weight_mem[16'h0944] <= 0;
        weight_mem[16'h0945] <= 0;
        weight_mem[16'h0946] <= 0;
        weight_mem[16'h0947] <= 0;
        weight_mem[16'h0948] <= 0;
        weight_mem[16'h0949] <= 0;
        weight_mem[16'h094A] <= 0;
        weight_mem[16'h094B] <= 0;
        weight_mem[16'h094C] <= 0;
        weight_mem[16'h094D] <= 0;
        weight_mem[16'h094E] <= 0;
        weight_mem[16'h094F] <= 0;
        weight_mem[16'h0950] <= 0;
        weight_mem[16'h0951] <= 0;
        weight_mem[16'h0952] <= 0;
        weight_mem[16'h0953] <= 0;
        weight_mem[16'h0954] <= 0;
        weight_mem[16'h0955] <= 0;
        weight_mem[16'h0956] <= 0;
        weight_mem[16'h0957] <= 0;
        weight_mem[16'h0958] <= 0;
        weight_mem[16'h0959] <= 0;
        weight_mem[16'h095A] <= 0;
        weight_mem[16'h095B] <= 0;
        weight_mem[16'h095C] <= 0;
        weight_mem[16'h095D] <= 0;
        weight_mem[16'h095E] <= 0;
        weight_mem[16'h095F] <= 0;
        weight_mem[16'h0960] <= 0;
        weight_mem[16'h0961] <= 0;
        weight_mem[16'h0962] <= 0;
        weight_mem[16'h0963] <= 0;
        weight_mem[16'h0964] <= 0;
        weight_mem[16'h0965] <= 0;
        weight_mem[16'h0966] <= 0;
        weight_mem[16'h0967] <= 0;
        weight_mem[16'h0968] <= 0;
        weight_mem[16'h0969] <= 0;
        weight_mem[16'h096A] <= 0;
        weight_mem[16'h096B] <= 0;
        weight_mem[16'h096C] <= 0;
        weight_mem[16'h096D] <= 0;
        weight_mem[16'h096E] <= 0;
        weight_mem[16'h096F] <= 0;
        weight_mem[16'h0970] <= 0;
        weight_mem[16'h0971] <= 0;
        weight_mem[16'h0972] <= 0;
        weight_mem[16'h0973] <= 0;
        weight_mem[16'h0974] <= 0;
        weight_mem[16'h0975] <= 0;
        weight_mem[16'h0976] <= 0;
        weight_mem[16'h0977] <= 0;
        weight_mem[16'h0978] <= 0;
        weight_mem[16'h0979] <= 0;
        weight_mem[16'h097A] <= 0;
        weight_mem[16'h097B] <= 0;
        weight_mem[16'h097C] <= 0;
        weight_mem[16'h097D] <= 0;
        weight_mem[16'h097E] <= 0;
        weight_mem[16'h097F] <= 0;
        weight_mem[16'h0980] <= 0;
        weight_mem[16'h0981] <= 0;
        weight_mem[16'h0982] <= 0;
        weight_mem[16'h0983] <= 0;
        weight_mem[16'h0984] <= 0;
        weight_mem[16'h0985] <= 0;
        weight_mem[16'h0986] <= 0;
        weight_mem[16'h0987] <= 0;
        weight_mem[16'h0988] <= 0;
        weight_mem[16'h0989] <= 0;
        weight_mem[16'h098A] <= 0;
        weight_mem[16'h098B] <= 0;
        weight_mem[16'h098C] <= 0;
        weight_mem[16'h098D] <= 0;
        weight_mem[16'h098E] <= 0;
        weight_mem[16'h098F] <= 0;
        weight_mem[16'h0990] <= 0;
        weight_mem[16'h0991] <= 0;
        weight_mem[16'h0992] <= 0;
        weight_mem[16'h0993] <= 0;
        weight_mem[16'h0994] <= 0;
        weight_mem[16'h0995] <= 0;
        weight_mem[16'h0996] <= 0;
        weight_mem[16'h0997] <= 0;
        weight_mem[16'h0998] <= 0;
        weight_mem[16'h0999] <= 0;
        weight_mem[16'h099A] <= 0;
        weight_mem[16'h099B] <= 0;
        weight_mem[16'h099C] <= 0;
        weight_mem[16'h099D] <= 0;
        weight_mem[16'h099E] <= 0;
        weight_mem[16'h099F] <= 0;
        weight_mem[16'h09A0] <= 0;
        weight_mem[16'h09A1] <= 0;
        weight_mem[16'h09A2] <= 0;
        weight_mem[16'h09A3] <= 0;
        weight_mem[16'h09A4] <= 0;
        weight_mem[16'h09A5] <= 0;
        weight_mem[16'h09A6] <= 0;
        weight_mem[16'h09A7] <= 0;
        weight_mem[16'h09A8] <= 0;
        weight_mem[16'h09A9] <= 0;
        weight_mem[16'h09AA] <= 0;
        weight_mem[16'h09AB] <= 0;
        weight_mem[16'h09AC] <= 0;
        weight_mem[16'h09AD] <= 0;
        weight_mem[16'h09AE] <= 0;
        weight_mem[16'h09AF] <= 0;

        // layer 1 neuron 5
        weight_mem[16'h0A00] <= 0;
        weight_mem[16'h0A01] <= 0;
        weight_mem[16'h0A02] <= 0;
        weight_mem[16'h0A03] <= 0;
        weight_mem[16'h0A04] <= 0;
        weight_mem[16'h0A05] <= 0;
        weight_mem[16'h0A06] <= 0;
        weight_mem[16'h0A07] <= 0;
        weight_mem[16'h0A08] <= 0;
        weight_mem[16'h0A09] <= 0;
        weight_mem[16'h0A0A] <= 0;
        weight_mem[16'h0A0B] <= 0;
        weight_mem[16'h0A0C] <= 0;
        weight_mem[16'h0A0D] <= 0;
        weight_mem[16'h0A0E] <= 0;
        weight_mem[16'h0A0F] <= 0;
        weight_mem[16'h0A10] <= 0;
        weight_mem[16'h0A11] <= 0;
        weight_mem[16'h0A12] <= 0;
        weight_mem[16'h0A13] <= 0;
        weight_mem[16'h0A14] <= 0;
        weight_mem[16'h0A15] <= 0;
        weight_mem[16'h0A16] <= 0;
        weight_mem[16'h0A17] <= 0;
        weight_mem[16'h0A18] <= 0;
        weight_mem[16'h0A19] <= 0;
        weight_mem[16'h0A1A] <= 0;
        weight_mem[16'h0A1B] <= 0;
        weight_mem[16'h0A1C] <= 0;
        weight_mem[16'h0A1D] <= 0;
        weight_mem[16'h0A1E] <= 0;
        weight_mem[16'h0A1F] <= 0;
        weight_mem[16'h0A20] <= 0;
        weight_mem[16'h0A21] <= 0;
        weight_mem[16'h0A22] <= 0;
        weight_mem[16'h0A23] <= 0;
        weight_mem[16'h0A24] <= 0;
        weight_mem[16'h0A25] <= 0;
        weight_mem[16'h0A26] <= 0;
        weight_mem[16'h0A27] <= 0;
        weight_mem[16'h0A28] <= 0;
        weight_mem[16'h0A29] <= 0;
        weight_mem[16'h0A2A] <= 0;
        weight_mem[16'h0A2B] <= 0;
        weight_mem[16'h0A2C] <= 0;
        weight_mem[16'h0A2D] <= 0;
        weight_mem[16'h0A2E] <= 0;
        weight_mem[16'h0A2F] <= 0;
        weight_mem[16'h0A30] <= 0;
        weight_mem[16'h0A31] <= 0;
        weight_mem[16'h0A32] <= 0;
        weight_mem[16'h0A33] <= 0;
        weight_mem[16'h0A34] <= 0;
        weight_mem[16'h0A35] <= 0;
        weight_mem[16'h0A36] <= 0;
        weight_mem[16'h0A37] <= 0;
        weight_mem[16'h0A38] <= 0;
        weight_mem[16'h0A39] <= 0;
        weight_mem[16'h0A3A] <= 0;
        weight_mem[16'h0A3B] <= 0;
        weight_mem[16'h0A3C] <= 0;
        weight_mem[16'h0A3D] <= 0;
        weight_mem[16'h0A3E] <= 0;
        weight_mem[16'h0A3F] <= 0;
        weight_mem[16'h0A40] <= 0;
        weight_mem[16'h0A41] <= 0;
        weight_mem[16'h0A42] <= 0;
        weight_mem[16'h0A43] <= 0;
        weight_mem[16'h0A44] <= 0;
        weight_mem[16'h0A45] <= 0;
        weight_mem[16'h0A46] <= 0;
        weight_mem[16'h0A47] <= 0;
        weight_mem[16'h0A48] <= 0;
        weight_mem[16'h0A49] <= 0;
        weight_mem[16'h0A4A] <= 0;
        weight_mem[16'h0A4B] <= 0;
        weight_mem[16'h0A4C] <= 0;
        weight_mem[16'h0A4D] <= 0;
        weight_mem[16'h0A4E] <= 0;
        weight_mem[16'h0A4F] <= 0;
        weight_mem[16'h0A50] <= 0;
        weight_mem[16'h0A51] <= 0;
        weight_mem[16'h0A52] <= 0;
        weight_mem[16'h0A53] <= 0;
        weight_mem[16'h0A54] <= 0;
        weight_mem[16'h0A55] <= 0;
        weight_mem[16'h0A56] <= 0;
        weight_mem[16'h0A57] <= 0;
        weight_mem[16'h0A58] <= 0;
        weight_mem[16'h0A59] <= 0;
        weight_mem[16'h0A5A] <= 0;
        weight_mem[16'h0A5B] <= 0;
        weight_mem[16'h0A5C] <= 0;
        weight_mem[16'h0A5D] <= 0;
        weight_mem[16'h0A5E] <= 0;
        weight_mem[16'h0A5F] <= 0;
        weight_mem[16'h0A60] <= 0;
        weight_mem[16'h0A61] <= 0;
        weight_mem[16'h0A62] <= 0;
        weight_mem[16'h0A63] <= 0;
        weight_mem[16'h0A64] <= 0;
        weight_mem[16'h0A65] <= 0;
        weight_mem[16'h0A66] <= 0;
        weight_mem[16'h0A67] <= 0;
        weight_mem[16'h0A68] <= 0;
        weight_mem[16'h0A69] <= 0;
        weight_mem[16'h0A6A] <= 0;
        weight_mem[16'h0A6B] <= 0;
        weight_mem[16'h0A6C] <= 0;
        weight_mem[16'h0A6D] <= 0;
        weight_mem[16'h0A6E] <= 0;
        weight_mem[16'h0A6F] <= 0;
        weight_mem[16'h0A70] <= 0;
        weight_mem[16'h0A71] <= 0;
        weight_mem[16'h0A72] <= 0;
        weight_mem[16'h0A73] <= 0;
        weight_mem[16'h0A74] <= 0;
        weight_mem[16'h0A75] <= 0;
        weight_mem[16'h0A76] <= 0;
        weight_mem[16'h0A77] <= 0;
        weight_mem[16'h0A78] <= 0;
        weight_mem[16'h0A79] <= 0;
        weight_mem[16'h0A7A] <= 0;
        weight_mem[16'h0A7B] <= 0;
        weight_mem[16'h0A7C] <= 0;
        weight_mem[16'h0A7D] <= 0;
        weight_mem[16'h0A7E] <= 0;
        weight_mem[16'h0A7F] <= 0;
        weight_mem[16'h0A80] <= 0;
        weight_mem[16'h0A81] <= 0;
        weight_mem[16'h0A82] <= 0;
        weight_mem[16'h0A83] <= 0;
        weight_mem[16'h0A84] <= 0;
        weight_mem[16'h0A85] <= 0;
        weight_mem[16'h0A86] <= 0;
        weight_mem[16'h0A87] <= 0;
        weight_mem[16'h0A88] <= 0;
        weight_mem[16'h0A89] <= 0;
        weight_mem[16'h0A8A] <= 0;
        weight_mem[16'h0A8B] <= 0;
        weight_mem[16'h0A8C] <= 0;
        weight_mem[16'h0A8D] <= 0;
        weight_mem[16'h0A8E] <= 0;
        weight_mem[16'h0A8F] <= 0;
        weight_mem[16'h0A90] <= 0;
        weight_mem[16'h0A91] <= 0;
        weight_mem[16'h0A92] <= 0;
        weight_mem[16'h0A93] <= 0;
        weight_mem[16'h0A94] <= 0;
        weight_mem[16'h0A95] <= 0;
        weight_mem[16'h0A96] <= 0;
        weight_mem[16'h0A97] <= 0;
        weight_mem[16'h0A98] <= 0;
        weight_mem[16'h0A99] <= 0;
        weight_mem[16'h0A9A] <= 0;
        weight_mem[16'h0A9B] <= 0;
        weight_mem[16'h0A9C] <= 0;
        weight_mem[16'h0A9D] <= 0;
        weight_mem[16'h0A9E] <= 0;
        weight_mem[16'h0A9F] <= 0;
        weight_mem[16'h0AA0] <= 0;
        weight_mem[16'h0AA1] <= 0;
        weight_mem[16'h0AA2] <= 0;
        weight_mem[16'h0AA3] <= 0;
        weight_mem[16'h0AA4] <= 0;
        weight_mem[16'h0AA5] <= 0;
        weight_mem[16'h0AA6] <= 0;
        weight_mem[16'h0AA7] <= 0;
        weight_mem[16'h0AA8] <= 0;
        weight_mem[16'h0AA9] <= 0;
        weight_mem[16'h0AAA] <= 0;
        weight_mem[16'h0AAB] <= 0;
        weight_mem[16'h0AAC] <= 0;
        weight_mem[16'h0AAD] <= 0;
        weight_mem[16'h0AAE] <= 0;
        weight_mem[16'h0AAF] <= 0;
        weight_mem[16'h0AB0] <= 0;
        weight_mem[16'h0AB1] <= 0;
        weight_mem[16'h0AB2] <= 0;
        weight_mem[16'h0AB3] <= 0;
        weight_mem[16'h0AB4] <= 0;
        weight_mem[16'h0AB5] <= 0;
        weight_mem[16'h0AB6] <= 0;
        weight_mem[16'h0AB7] <= 0;
        weight_mem[16'h0AB8] <= 0;
        weight_mem[16'h0AB9] <= 0;
        weight_mem[16'h0ABA] <= 0;
        weight_mem[16'h0ABB] <= 0;
        weight_mem[16'h0ABC] <= 0;
        weight_mem[16'h0ABD] <= 0;
        weight_mem[16'h0ABE] <= 0;
        weight_mem[16'h0ABF] <= 0;
        weight_mem[16'h0AC0] <= 0;
        weight_mem[16'h0AC1] <= 0;
        weight_mem[16'h0AC2] <= 0;
        weight_mem[16'h0AC3] <= 0;
        weight_mem[16'h0AC4] <= 0;
        weight_mem[16'h0AC5] <= 0;
        weight_mem[16'h0AC6] <= 0;
        weight_mem[16'h0AC7] <= 0;
        weight_mem[16'h0AC8] <= 0;
        weight_mem[16'h0AC9] <= 0;
        weight_mem[16'h0ACA] <= 0;
        weight_mem[16'h0ACB] <= 0;
        weight_mem[16'h0ACC] <= 0;
        weight_mem[16'h0ACD] <= 0;
        weight_mem[16'h0ACE] <= 0;
        weight_mem[16'h0ACF] <= 0;
        weight_mem[16'h0AD0] <= 0;
        weight_mem[16'h0AD1] <= 0;
        weight_mem[16'h0AD2] <= 0;
        weight_mem[16'h0AD3] <= 0;
        weight_mem[16'h0AD4] <= 0;
        weight_mem[16'h0AD5] <= 0;
        weight_mem[16'h0AD6] <= 0;
        weight_mem[16'h0AD7] <= 0;
        weight_mem[16'h0AD8] <= 0;
        weight_mem[16'h0AD9] <= 0;
        weight_mem[16'h0ADA] <= 0;
        weight_mem[16'h0ADB] <= 0;
        weight_mem[16'h0ADC] <= 0;
        weight_mem[16'h0ADD] <= 0;
        weight_mem[16'h0ADE] <= 0;
        weight_mem[16'h0ADF] <= 0;
        weight_mem[16'h0AE0] <= 0;
        weight_mem[16'h0AE1] <= 0;
        weight_mem[16'h0AE2] <= 0;
        weight_mem[16'h0AE3] <= 0;
        weight_mem[16'h0AE4] <= 0;
        weight_mem[16'h0AE5] <= 0;
        weight_mem[16'h0AE6] <= 0;
        weight_mem[16'h0AE7] <= 0;
        weight_mem[16'h0AE8] <= 0;
        weight_mem[16'h0AE9] <= 0;
        weight_mem[16'h0AEA] <= 0;
        weight_mem[16'h0AEB] <= 0;
        weight_mem[16'h0AEC] <= 0;
        weight_mem[16'h0AED] <= 0;
        weight_mem[16'h0AEE] <= 0;
        weight_mem[16'h0AEF] <= 0;
        weight_mem[16'h0AF0] <= 0;
        weight_mem[16'h0AF1] <= 0;
        weight_mem[16'h0AF2] <= 0;
        weight_mem[16'h0AF3] <= 0;
        weight_mem[16'h0AF4] <= 0;
        weight_mem[16'h0AF5] <= 0;
        weight_mem[16'h0AF6] <= 0;
        weight_mem[16'h0AF7] <= 0;
        weight_mem[16'h0AF8] <= 0;
        weight_mem[16'h0AF9] <= 0;
        weight_mem[16'h0AFA] <= 0;
        weight_mem[16'h0AFB] <= 0;
        weight_mem[16'h0AFC] <= 0;
        weight_mem[16'h0AFD] <= 0;
        weight_mem[16'h0AFE] <= 0;
        weight_mem[16'h0AFF] <= 0;
        weight_mem[16'h0B00] <= 0;
        weight_mem[16'h0B01] <= 0;
        weight_mem[16'h0B02] <= 0;
        weight_mem[16'h0B03] <= 0;
        weight_mem[16'h0B04] <= 0;
        weight_mem[16'h0B05] <= 0;
        weight_mem[16'h0B06] <= 0;
        weight_mem[16'h0B07] <= 0;
        weight_mem[16'h0B08] <= 0;
        weight_mem[16'h0B09] <= 0;
        weight_mem[16'h0B0A] <= 0;
        weight_mem[16'h0B0B] <= 0;
        weight_mem[16'h0B0C] <= 0;
        weight_mem[16'h0B0D] <= 0;
        weight_mem[16'h0B0E] <= 0;
        weight_mem[16'h0B0F] <= 0;
        weight_mem[16'h0B10] <= 0;
        weight_mem[16'h0B11] <= 0;
        weight_mem[16'h0B12] <= 0;
        weight_mem[16'h0B13] <= 0;
        weight_mem[16'h0B14] <= 0;
        weight_mem[16'h0B15] <= 0;
        weight_mem[16'h0B16] <= 0;
        weight_mem[16'h0B17] <= 0;
        weight_mem[16'h0B18] <= 0;
        weight_mem[16'h0B19] <= 0;
        weight_mem[16'h0B1A] <= 0;
        weight_mem[16'h0B1B] <= 0;
        weight_mem[16'h0B1C] <= 0;
        weight_mem[16'h0B1D] <= 0;
        weight_mem[16'h0B1E] <= 0;
        weight_mem[16'h0B1F] <= 0;
        weight_mem[16'h0B20] <= 0;
        weight_mem[16'h0B21] <= 0;
        weight_mem[16'h0B22] <= 0;
        weight_mem[16'h0B23] <= 0;
        weight_mem[16'h0B24] <= 0;
        weight_mem[16'h0B25] <= 0;
        weight_mem[16'h0B26] <= 0;
        weight_mem[16'h0B27] <= 0;
        weight_mem[16'h0B28] <= 0;
        weight_mem[16'h0B29] <= 0;
        weight_mem[16'h0B2A] <= 0;
        weight_mem[16'h0B2B] <= 0;
        weight_mem[16'h0B2C] <= 0;
        weight_mem[16'h0B2D] <= 0;
        weight_mem[16'h0B2E] <= 0;
        weight_mem[16'h0B2F] <= 0;
        weight_mem[16'h0B30] <= 0;
        weight_mem[16'h0B31] <= 0;
        weight_mem[16'h0B32] <= 0;
        weight_mem[16'h0B33] <= 0;
        weight_mem[16'h0B34] <= 0;
        weight_mem[16'h0B35] <= 0;
        weight_mem[16'h0B36] <= 0;
        weight_mem[16'h0B37] <= 0;
        weight_mem[16'h0B38] <= 0;
        weight_mem[16'h0B39] <= 0;
        weight_mem[16'h0B3A] <= 0;
        weight_mem[16'h0B3B] <= 0;
        weight_mem[16'h0B3C] <= 0;
        weight_mem[16'h0B3D] <= 0;
        weight_mem[16'h0B3E] <= 0;
        weight_mem[16'h0B3F] <= 0;
        weight_mem[16'h0B40] <= 0;
        weight_mem[16'h0B41] <= 0;
        weight_mem[16'h0B42] <= 0;
        weight_mem[16'h0B43] <= 0;
        weight_mem[16'h0B44] <= 0;
        weight_mem[16'h0B45] <= 0;
        weight_mem[16'h0B46] <= 0;
        weight_mem[16'h0B47] <= 0;
        weight_mem[16'h0B48] <= 0;
        weight_mem[16'h0B49] <= 0;
        weight_mem[16'h0B4A] <= 0;
        weight_mem[16'h0B4B] <= 0;
        weight_mem[16'h0B4C] <= 0;
        weight_mem[16'h0B4D] <= 0;
        weight_mem[16'h0B4E] <= 0;
        weight_mem[16'h0B4F] <= 0;
        weight_mem[16'h0B50] <= 0;
        weight_mem[16'h0B51] <= 0;
        weight_mem[16'h0B52] <= 0;
        weight_mem[16'h0B53] <= 0;
        weight_mem[16'h0B54] <= 0;
        weight_mem[16'h0B55] <= 0;
        weight_mem[16'h0B56] <= 0;
        weight_mem[16'h0B57] <= 0;
        weight_mem[16'h0B58] <= 0;
        weight_mem[16'h0B59] <= 0;
        weight_mem[16'h0B5A] <= 0;
        weight_mem[16'h0B5B] <= 0;
        weight_mem[16'h0B5C] <= 0;
        weight_mem[16'h0B5D] <= 0;
        weight_mem[16'h0B5E] <= 0;
        weight_mem[16'h0B5F] <= 0;
        weight_mem[16'h0B60] <= 0;
        weight_mem[16'h0B61] <= 0;
        weight_mem[16'h0B62] <= 0;
        weight_mem[16'h0B63] <= 0;
        weight_mem[16'h0B64] <= 0;
        weight_mem[16'h0B65] <= 0;
        weight_mem[16'h0B66] <= 0;
        weight_mem[16'h0B67] <= 0;
        weight_mem[16'h0B68] <= 0;
        weight_mem[16'h0B69] <= 0;
        weight_mem[16'h0B6A] <= 0;
        weight_mem[16'h0B6B] <= 0;
        weight_mem[16'h0B6C] <= 0;
        weight_mem[16'h0B6D] <= 0;
        weight_mem[16'h0B6E] <= 0;
        weight_mem[16'h0B6F] <= 0;
        weight_mem[16'h0B70] <= 0;
        weight_mem[16'h0B71] <= 0;
        weight_mem[16'h0B72] <= 0;
        weight_mem[16'h0B73] <= 0;
        weight_mem[16'h0B74] <= 0;
        weight_mem[16'h0B75] <= 0;
        weight_mem[16'h0B76] <= 0;
        weight_mem[16'h0B77] <= 0;
        weight_mem[16'h0B78] <= 0;
        weight_mem[16'h0B79] <= 0;
        weight_mem[16'h0B7A] <= 0;
        weight_mem[16'h0B7B] <= 0;
        weight_mem[16'h0B7C] <= 0;
        weight_mem[16'h0B7D] <= 0;
        weight_mem[16'h0B7E] <= 0;
        weight_mem[16'h0B7F] <= 0;
        weight_mem[16'h0B80] <= 0;
        weight_mem[16'h0B81] <= 0;
        weight_mem[16'h0B82] <= 0;
        weight_mem[16'h0B83] <= 0;
        weight_mem[16'h0B84] <= 0;
        weight_mem[16'h0B85] <= 0;
        weight_mem[16'h0B86] <= 0;
        weight_mem[16'h0B87] <= 0;
        weight_mem[16'h0B88] <= 0;
        weight_mem[16'h0B89] <= 0;
        weight_mem[16'h0B8A] <= 0;
        weight_mem[16'h0B8B] <= 0;
        weight_mem[16'h0B8C] <= 0;
        weight_mem[16'h0B8D] <= 0;
        weight_mem[16'h0B8E] <= 0;
        weight_mem[16'h0B8F] <= 0;
        weight_mem[16'h0B90] <= 0;
        weight_mem[16'h0B91] <= 0;
        weight_mem[16'h0B92] <= 0;
        weight_mem[16'h0B93] <= 0;
        weight_mem[16'h0B94] <= 0;
        weight_mem[16'h0B95] <= 0;
        weight_mem[16'h0B96] <= 0;
        weight_mem[16'h0B97] <= 0;
        weight_mem[16'h0B98] <= 0;
        weight_mem[16'h0B99] <= 0;
        weight_mem[16'h0B9A] <= 0;
        weight_mem[16'h0B9B] <= 0;
        weight_mem[16'h0B9C] <= 0;
        weight_mem[16'h0B9D] <= 0;
        weight_mem[16'h0B9E] <= 0;
        weight_mem[16'h0B9F] <= 0;
        weight_mem[16'h0BA0] <= 0;
        weight_mem[16'h0BA1] <= 0;
        weight_mem[16'h0BA2] <= 0;
        weight_mem[16'h0BA3] <= 0;
        weight_mem[16'h0BA4] <= 0;
        weight_mem[16'h0BA5] <= 0;
        weight_mem[16'h0BA6] <= 0;
        weight_mem[16'h0BA7] <= 0;
        weight_mem[16'h0BA8] <= 0;
        weight_mem[16'h0BA9] <= 0;
        weight_mem[16'h0BAA] <= 0;
        weight_mem[16'h0BAB] <= 0;
        weight_mem[16'h0BAC] <= 0;
        weight_mem[16'h0BAD] <= 0;
        weight_mem[16'h0BAE] <= 0;
        weight_mem[16'h0BAF] <= 0;

        // layer 1 neuron 6
        weight_mem[16'h0C00] <= 0;
        weight_mem[16'h0C01] <= 0;
        weight_mem[16'h0C02] <= 0;
        weight_mem[16'h0C03] <= 0;
        weight_mem[16'h0C04] <= 0;
        weight_mem[16'h0C05] <= 0;
        weight_mem[16'h0C06] <= 0;
        weight_mem[16'h0C07] <= 0;
        weight_mem[16'h0C08] <= 0;
        weight_mem[16'h0C09] <= 0;
        weight_mem[16'h0C0A] <= 0;
        weight_mem[16'h0C0B] <= 0;
        weight_mem[16'h0C0C] <= 0;
        weight_mem[16'h0C0D] <= 0;
        weight_mem[16'h0C0E] <= 0;
        weight_mem[16'h0C0F] <= 0;
        weight_mem[16'h0C10] <= 0;
        weight_mem[16'h0C11] <= 0;
        weight_mem[16'h0C12] <= 0;
        weight_mem[16'h0C13] <= 0;
        weight_mem[16'h0C14] <= 0;
        weight_mem[16'h0C15] <= 0;
        weight_mem[16'h0C16] <= 0;
        weight_mem[16'h0C17] <= 0;
        weight_mem[16'h0C18] <= 0;
        weight_mem[16'h0C19] <= 0;
        weight_mem[16'h0C1A] <= 0;
        weight_mem[16'h0C1B] <= 0;
        weight_mem[16'h0C1C] <= 0;
        weight_mem[16'h0C1D] <= 0;
        weight_mem[16'h0C1E] <= 0;
        weight_mem[16'h0C1F] <= 0;
        weight_mem[16'h0C20] <= 0;
        weight_mem[16'h0C21] <= 0;
        weight_mem[16'h0C22] <= 0;
        weight_mem[16'h0C23] <= 0;
        weight_mem[16'h0C24] <= 0;
        weight_mem[16'h0C25] <= 0;
        weight_mem[16'h0C26] <= 0;
        weight_mem[16'h0C27] <= 0;
        weight_mem[16'h0C28] <= 0;
        weight_mem[16'h0C29] <= 0;
        weight_mem[16'h0C2A] <= 0;
        weight_mem[16'h0C2B] <= 0;
        weight_mem[16'h0C2C] <= 0;
        weight_mem[16'h0C2D] <= 0;
        weight_mem[16'h0C2E] <= 0;
        weight_mem[16'h0C2F] <= 0;
        weight_mem[16'h0C30] <= 0;
        weight_mem[16'h0C31] <= 0;
        weight_mem[16'h0C32] <= 0;
        weight_mem[16'h0C33] <= 0;
        weight_mem[16'h0C34] <= 0;
        weight_mem[16'h0C35] <= 0;
        weight_mem[16'h0C36] <= 0;
        weight_mem[16'h0C37] <= 0;
        weight_mem[16'h0C38] <= 0;
        weight_mem[16'h0C39] <= 0;
        weight_mem[16'h0C3A] <= 0;
        weight_mem[16'h0C3B] <= 0;
        weight_mem[16'h0C3C] <= 0;
        weight_mem[16'h0C3D] <= 0;
        weight_mem[16'h0C3E] <= 0;
        weight_mem[16'h0C3F] <= 0;
        weight_mem[16'h0C40] <= 0;
        weight_mem[16'h0C41] <= 0;
        weight_mem[16'h0C42] <= 0;
        weight_mem[16'h0C43] <= 0;
        weight_mem[16'h0C44] <= 0;
        weight_mem[16'h0C45] <= 0;
        weight_mem[16'h0C46] <= 0;
        weight_mem[16'h0C47] <= 0;
        weight_mem[16'h0C48] <= 0;
        weight_mem[16'h0C49] <= 0;
        weight_mem[16'h0C4A] <= 0;
        weight_mem[16'h0C4B] <= 0;
        weight_mem[16'h0C4C] <= 0;
        weight_mem[16'h0C4D] <= 0;
        weight_mem[16'h0C4E] <= 0;
        weight_mem[16'h0C4F] <= 0;
        weight_mem[16'h0C50] <= 0;
        weight_mem[16'h0C51] <= 0;
        weight_mem[16'h0C52] <= 0;
        weight_mem[16'h0C53] <= 0;
        weight_mem[16'h0C54] <= 0;
        weight_mem[16'h0C55] <= 0;
        weight_mem[16'h0C56] <= 0;
        weight_mem[16'h0C57] <= 0;
        weight_mem[16'h0C58] <= 0;
        weight_mem[16'h0C59] <= 0;
        weight_mem[16'h0C5A] <= 0;
        weight_mem[16'h0C5B] <= 0;
        weight_mem[16'h0C5C] <= 0;
        weight_mem[16'h0C5D] <= 0;
        weight_mem[16'h0C5E] <= 0;
        weight_mem[16'h0C5F] <= 0;
        weight_mem[16'h0C60] <= 0;
        weight_mem[16'h0C61] <= 0;
        weight_mem[16'h0C62] <= 0;
        weight_mem[16'h0C63] <= 0;
        weight_mem[16'h0C64] <= 0;
        weight_mem[16'h0C65] <= 0;
        weight_mem[16'h0C66] <= 0;
        weight_mem[16'h0C67] <= 0;
        weight_mem[16'h0C68] <= 0;
        weight_mem[16'h0C69] <= 0;
        weight_mem[16'h0C6A] <= 0;
        weight_mem[16'h0C6B] <= 0;
        weight_mem[16'h0C6C] <= 0;
        weight_mem[16'h0C6D] <= 0;
        weight_mem[16'h0C6E] <= 0;
        weight_mem[16'h0C6F] <= 0;
        weight_mem[16'h0C70] <= 0;
        weight_mem[16'h0C71] <= 0;
        weight_mem[16'h0C72] <= 0;
        weight_mem[16'h0C73] <= 0;
        weight_mem[16'h0C74] <= 0;
        weight_mem[16'h0C75] <= 0;
        weight_mem[16'h0C76] <= 0;
        weight_mem[16'h0C77] <= 0;
        weight_mem[16'h0C78] <= 0;
        weight_mem[16'h0C79] <= 0;
        weight_mem[16'h0C7A] <= 0;
        weight_mem[16'h0C7B] <= 0;
        weight_mem[16'h0C7C] <= 0;
        weight_mem[16'h0C7D] <= 0;
        weight_mem[16'h0C7E] <= 0;
        weight_mem[16'h0C7F] <= 0;
        weight_mem[16'h0C80] <= 0;
        weight_mem[16'h0C81] <= 0;
        weight_mem[16'h0C82] <= 0;
        weight_mem[16'h0C83] <= 0;
        weight_mem[16'h0C84] <= 0;
        weight_mem[16'h0C85] <= 0;
        weight_mem[16'h0C86] <= 0;
        weight_mem[16'h0C87] <= 0;
        weight_mem[16'h0C88] <= 0;
        weight_mem[16'h0C89] <= 0;
        weight_mem[16'h0C8A] <= 0;
        weight_mem[16'h0C8B] <= 0;
        weight_mem[16'h0C8C] <= 0;
        weight_mem[16'h0C8D] <= 0;
        weight_mem[16'h0C8E] <= 0;
        weight_mem[16'h0C8F] <= 0;
        weight_mem[16'h0C90] <= 0;
        weight_mem[16'h0C91] <= 0;
        weight_mem[16'h0C92] <= 0;
        weight_mem[16'h0C93] <= 0;
        weight_mem[16'h0C94] <= 0;
        weight_mem[16'h0C95] <= 0;
        weight_mem[16'h0C96] <= 0;
        weight_mem[16'h0C97] <= 0;
        weight_mem[16'h0C98] <= 0;
        weight_mem[16'h0C99] <= 0;
        weight_mem[16'h0C9A] <= 0;
        weight_mem[16'h0C9B] <= 0;
        weight_mem[16'h0C9C] <= 0;
        weight_mem[16'h0C9D] <= 0;
        weight_mem[16'h0C9E] <= 0;
        weight_mem[16'h0C9F] <= 0;
        weight_mem[16'h0CA0] <= 0;
        weight_mem[16'h0CA1] <= 0;
        weight_mem[16'h0CA2] <= 0;
        weight_mem[16'h0CA3] <= 0;
        weight_mem[16'h0CA4] <= 0;
        weight_mem[16'h0CA5] <= 0;
        weight_mem[16'h0CA6] <= 0;
        weight_mem[16'h0CA7] <= 0;
        weight_mem[16'h0CA8] <= 0;
        weight_mem[16'h0CA9] <= 0;
        weight_mem[16'h0CAA] <= 0;
        weight_mem[16'h0CAB] <= 0;
        weight_mem[16'h0CAC] <= 0;
        weight_mem[16'h0CAD] <= 0;
        weight_mem[16'h0CAE] <= 0;
        weight_mem[16'h0CAF] <= 0;
        weight_mem[16'h0CB0] <= 0;
        weight_mem[16'h0CB1] <= 0;
        weight_mem[16'h0CB2] <= 0;
        weight_mem[16'h0CB3] <= 0;
        weight_mem[16'h0CB4] <= 0;
        weight_mem[16'h0CB5] <= 0;
        weight_mem[16'h0CB6] <= 0;
        weight_mem[16'h0CB7] <= 0;
        weight_mem[16'h0CB8] <= 0;
        weight_mem[16'h0CB9] <= 0;
        weight_mem[16'h0CBA] <= 0;
        weight_mem[16'h0CBB] <= 0;
        weight_mem[16'h0CBC] <= 0;
        weight_mem[16'h0CBD] <= 0;
        weight_mem[16'h0CBE] <= 0;
        weight_mem[16'h0CBF] <= 0;
        weight_mem[16'h0CC0] <= 0;
        weight_mem[16'h0CC1] <= 0;
        weight_mem[16'h0CC2] <= 0;
        weight_mem[16'h0CC3] <= 0;
        weight_mem[16'h0CC4] <= 0;
        weight_mem[16'h0CC5] <= 0;
        weight_mem[16'h0CC6] <= 0;
        weight_mem[16'h0CC7] <= 0;
        weight_mem[16'h0CC8] <= 0;
        weight_mem[16'h0CC9] <= 0;
        weight_mem[16'h0CCA] <= 0;
        weight_mem[16'h0CCB] <= 0;
        weight_mem[16'h0CCC] <= 0;
        weight_mem[16'h0CCD] <= 0;
        weight_mem[16'h0CCE] <= 0;
        weight_mem[16'h0CCF] <= 0;
        weight_mem[16'h0CD0] <= 0;
        weight_mem[16'h0CD1] <= 0;
        weight_mem[16'h0CD2] <= 0;
        weight_mem[16'h0CD3] <= 0;
        weight_mem[16'h0CD4] <= 0;
        weight_mem[16'h0CD5] <= 0;
        weight_mem[16'h0CD6] <= 0;
        weight_mem[16'h0CD7] <= 0;
        weight_mem[16'h0CD8] <= 0;
        weight_mem[16'h0CD9] <= 0;
        weight_mem[16'h0CDA] <= 0;
        weight_mem[16'h0CDB] <= 0;
        weight_mem[16'h0CDC] <= 0;
        weight_mem[16'h0CDD] <= 0;
        weight_mem[16'h0CDE] <= 0;
        weight_mem[16'h0CDF] <= 0;
        weight_mem[16'h0CE0] <= 0;
        weight_mem[16'h0CE1] <= 0;
        weight_mem[16'h0CE2] <= 0;
        weight_mem[16'h0CE3] <= 0;
        weight_mem[16'h0CE4] <= 0;
        weight_mem[16'h0CE5] <= 0;
        weight_mem[16'h0CE6] <= 0;
        weight_mem[16'h0CE7] <= 0;
        weight_mem[16'h0CE8] <= 0;
        weight_mem[16'h0CE9] <= 0;
        weight_mem[16'h0CEA] <= 0;
        weight_mem[16'h0CEB] <= 0;
        weight_mem[16'h0CEC] <= 0;
        weight_mem[16'h0CED] <= 0;
        weight_mem[16'h0CEE] <= 0;
        weight_mem[16'h0CEF] <= 0;
        weight_mem[16'h0CF0] <= 0;
        weight_mem[16'h0CF1] <= 0;
        weight_mem[16'h0CF2] <= 0;
        weight_mem[16'h0CF3] <= 0;
        weight_mem[16'h0CF4] <= 0;
        weight_mem[16'h0CF5] <= 0;
        weight_mem[16'h0CF6] <= 0;
        weight_mem[16'h0CF7] <= 0;
        weight_mem[16'h0CF8] <= 0;
        weight_mem[16'h0CF9] <= 0;
        weight_mem[16'h0CFA] <= 0;
        weight_mem[16'h0CFB] <= 0;
        weight_mem[16'h0CFC] <= 0;
        weight_mem[16'h0CFD] <= 0;
        weight_mem[16'h0CFE] <= 0;
        weight_mem[16'h0CFF] <= 0;
        weight_mem[16'h0D00] <= 0;
        weight_mem[16'h0D01] <= 0;
        weight_mem[16'h0D02] <= 0;
        weight_mem[16'h0D03] <= 0;
        weight_mem[16'h0D04] <= 0;
        weight_mem[16'h0D05] <= 0;
        weight_mem[16'h0D06] <= 0;
        weight_mem[16'h0D07] <= 0;
        weight_mem[16'h0D08] <= 0;
        weight_mem[16'h0D09] <= 0;
        weight_mem[16'h0D0A] <= 0;
        weight_mem[16'h0D0B] <= 0;
        weight_mem[16'h0D0C] <= 0;
        weight_mem[16'h0D0D] <= 0;
        weight_mem[16'h0D0E] <= 0;
        weight_mem[16'h0D0F] <= 0;
        weight_mem[16'h0D10] <= 0;
        weight_mem[16'h0D11] <= 0;
        weight_mem[16'h0D12] <= 0;
        weight_mem[16'h0D13] <= 0;
        weight_mem[16'h0D14] <= 0;
        weight_mem[16'h0D15] <= 0;
        weight_mem[16'h0D16] <= 0;
        weight_mem[16'h0D17] <= 0;
        weight_mem[16'h0D18] <= 0;
        weight_mem[16'h0D19] <= 0;
        weight_mem[16'h0D1A] <= 0;
        weight_mem[16'h0D1B] <= 0;
        weight_mem[16'h0D1C] <= 0;
        weight_mem[16'h0D1D] <= 0;
        weight_mem[16'h0D1E] <= 0;
        weight_mem[16'h0D1F] <= 0;
        weight_mem[16'h0D20] <= 0;
        weight_mem[16'h0D21] <= 0;
        weight_mem[16'h0D22] <= 0;
        weight_mem[16'h0D23] <= 0;
        weight_mem[16'h0D24] <= 0;
        weight_mem[16'h0D25] <= 0;
        weight_mem[16'h0D26] <= 0;
        weight_mem[16'h0D27] <= 0;
        weight_mem[16'h0D28] <= 0;
        weight_mem[16'h0D29] <= 0;
        weight_mem[16'h0D2A] <= 0;
        weight_mem[16'h0D2B] <= 0;
        weight_mem[16'h0D2C] <= 0;
        weight_mem[16'h0D2D] <= 0;
        weight_mem[16'h0D2E] <= 0;
        weight_mem[16'h0D2F] <= 0;
        weight_mem[16'h0D30] <= 0;
        weight_mem[16'h0D31] <= 0;
        weight_mem[16'h0D32] <= 0;
        weight_mem[16'h0D33] <= 0;
        weight_mem[16'h0D34] <= 0;
        weight_mem[16'h0D35] <= 0;
        weight_mem[16'h0D36] <= 0;
        weight_mem[16'h0D37] <= 0;
        weight_mem[16'h0D38] <= 0;
        weight_mem[16'h0D39] <= 0;
        weight_mem[16'h0D3A] <= 0;
        weight_mem[16'h0D3B] <= 0;
        weight_mem[16'h0D3C] <= 0;
        weight_mem[16'h0D3D] <= 0;
        weight_mem[16'h0D3E] <= 0;
        weight_mem[16'h0D3F] <= 0;
        weight_mem[16'h0D40] <= 0;
        weight_mem[16'h0D41] <= 0;
        weight_mem[16'h0D42] <= 0;
        weight_mem[16'h0D43] <= 0;
        weight_mem[16'h0D44] <= 0;
        weight_mem[16'h0D45] <= 0;
        weight_mem[16'h0D46] <= 0;
        weight_mem[16'h0D47] <= 0;
        weight_mem[16'h0D48] <= 0;
        weight_mem[16'h0D49] <= 0;
        weight_mem[16'h0D4A] <= 0;
        weight_mem[16'h0D4B] <= 0;
        weight_mem[16'h0D4C] <= 0;
        weight_mem[16'h0D4D] <= 0;
        weight_mem[16'h0D4E] <= 0;
        weight_mem[16'h0D4F] <= 0;
        weight_mem[16'h0D50] <= 0;
        weight_mem[16'h0D51] <= 0;
        weight_mem[16'h0D52] <= 0;
        weight_mem[16'h0D53] <= 0;
        weight_mem[16'h0D54] <= 0;
        weight_mem[16'h0D55] <= 0;
        weight_mem[16'h0D56] <= 0;
        weight_mem[16'h0D57] <= 0;
        weight_mem[16'h0D58] <= 0;
        weight_mem[16'h0D59] <= 0;
        weight_mem[16'h0D5A] <= 0;
        weight_mem[16'h0D5B] <= 0;
        weight_mem[16'h0D5C] <= 0;
        weight_mem[16'h0D5D] <= 0;
        weight_mem[16'h0D5E] <= 0;
        weight_mem[16'h0D5F] <= 0;
        weight_mem[16'h0D60] <= 0;
        weight_mem[16'h0D61] <= 0;
        weight_mem[16'h0D62] <= 0;
        weight_mem[16'h0D63] <= 0;
        weight_mem[16'h0D64] <= 0;
        weight_mem[16'h0D65] <= 0;
        weight_mem[16'h0D66] <= 0;
        weight_mem[16'h0D67] <= 0;
        weight_mem[16'h0D68] <= 0;
        weight_mem[16'h0D69] <= 0;
        weight_mem[16'h0D6A] <= 0;
        weight_mem[16'h0D6B] <= 0;
        weight_mem[16'h0D6C] <= 0;
        weight_mem[16'h0D6D] <= 0;
        weight_mem[16'h0D6E] <= 0;
        weight_mem[16'h0D6F] <= 0;
        weight_mem[16'h0D70] <= 0;
        weight_mem[16'h0D71] <= 0;
        weight_mem[16'h0D72] <= 0;
        weight_mem[16'h0D73] <= 0;
        weight_mem[16'h0D74] <= 0;
        weight_mem[16'h0D75] <= 0;
        weight_mem[16'h0D76] <= 0;
        weight_mem[16'h0D77] <= 0;
        weight_mem[16'h0D78] <= 0;
        weight_mem[16'h0D79] <= 0;
        weight_mem[16'h0D7A] <= 0;
        weight_mem[16'h0D7B] <= 0;
        weight_mem[16'h0D7C] <= 0;
        weight_mem[16'h0D7D] <= 0;
        weight_mem[16'h0D7E] <= 0;
        weight_mem[16'h0D7F] <= 0;
        weight_mem[16'h0D80] <= 0;
        weight_mem[16'h0D81] <= 0;
        weight_mem[16'h0D82] <= 0;
        weight_mem[16'h0D83] <= 0;
        weight_mem[16'h0D84] <= 0;
        weight_mem[16'h0D85] <= 0;
        weight_mem[16'h0D86] <= 0;
        weight_mem[16'h0D87] <= 0;
        weight_mem[16'h0D88] <= 0;
        weight_mem[16'h0D89] <= 0;
        weight_mem[16'h0D8A] <= 0;
        weight_mem[16'h0D8B] <= 0;
        weight_mem[16'h0D8C] <= 0;
        weight_mem[16'h0D8D] <= 0;
        weight_mem[16'h0D8E] <= 0;
        weight_mem[16'h0D8F] <= 0;
        weight_mem[16'h0D90] <= 0;
        weight_mem[16'h0D91] <= 0;
        weight_mem[16'h0D92] <= 0;
        weight_mem[16'h0D93] <= 0;
        weight_mem[16'h0D94] <= 0;
        weight_mem[16'h0D95] <= 0;
        weight_mem[16'h0D96] <= 0;
        weight_mem[16'h0D97] <= 0;
        weight_mem[16'h0D98] <= 0;
        weight_mem[16'h0D99] <= 0;
        weight_mem[16'h0D9A] <= 0;
        weight_mem[16'h0D9B] <= 0;
        weight_mem[16'h0D9C] <= 0;
        weight_mem[16'h0D9D] <= 0;
        weight_mem[16'h0D9E] <= 0;
        weight_mem[16'h0D9F] <= 0;
        weight_mem[16'h0DA0] <= 0;
        weight_mem[16'h0DA1] <= 0;
        weight_mem[16'h0DA2] <= 0;
        weight_mem[16'h0DA3] <= 0;
        weight_mem[16'h0DA4] <= 0;
        weight_mem[16'h0DA5] <= 0;
        weight_mem[16'h0DA6] <= 0;
        weight_mem[16'h0DA7] <= 0;
        weight_mem[16'h0DA8] <= 0;
        weight_mem[16'h0DA9] <= 0;
        weight_mem[16'h0DAA] <= 0;
        weight_mem[16'h0DAB] <= 0;
        weight_mem[16'h0DAC] <= 0;
        weight_mem[16'h0DAD] <= 0;
        weight_mem[16'h0DAE] <= 0;
        weight_mem[16'h0DAF] <= 0;

        // layer 1 neuron 7
        weight_mem[16'h0E00] <= 0;
        weight_mem[16'h0E01] <= 0;
        weight_mem[16'h0E02] <= 0;
        weight_mem[16'h0E03] <= 0;
        weight_mem[16'h0E04] <= 0;
        weight_mem[16'h0E05] <= 0;
        weight_mem[16'h0E06] <= 0;
        weight_mem[16'h0E07] <= 0;
        weight_mem[16'h0E08] <= 0;
        weight_mem[16'h0E09] <= 0;
        weight_mem[16'h0E0A] <= 0;
        weight_mem[16'h0E0B] <= 0;
        weight_mem[16'h0E0C] <= 0;
        weight_mem[16'h0E0D] <= 0;
        weight_mem[16'h0E0E] <= 0;
        weight_mem[16'h0E0F] <= 0;
        weight_mem[16'h0E10] <= 0;
        weight_mem[16'h0E11] <= 0;
        weight_mem[16'h0E12] <= 0;
        weight_mem[16'h0E13] <= 0;
        weight_mem[16'h0E14] <= 0;
        weight_mem[16'h0E15] <= 0;
        weight_mem[16'h0E16] <= 0;
        weight_mem[16'h0E17] <= 0;
        weight_mem[16'h0E18] <= 0;
        weight_mem[16'h0E19] <= 0;
        weight_mem[16'h0E1A] <= 0;
        weight_mem[16'h0E1B] <= 0;
        weight_mem[16'h0E1C] <= 0;
        weight_mem[16'h0E1D] <= 0;
        weight_mem[16'h0E1E] <= 0;
        weight_mem[16'h0E1F] <= 0;
        weight_mem[16'h0E20] <= 0;
        weight_mem[16'h0E21] <= 0;
        weight_mem[16'h0E22] <= 0;
        weight_mem[16'h0E23] <= 0;
        weight_mem[16'h0E24] <= 0;
        weight_mem[16'h0E25] <= 0;
        weight_mem[16'h0E26] <= 0;
        weight_mem[16'h0E27] <= 0;
        weight_mem[16'h0E28] <= 0;
        weight_mem[16'h0E29] <= 0;
        weight_mem[16'h0E2A] <= 0;
        weight_mem[16'h0E2B] <= 0;
        weight_mem[16'h0E2C] <= 0;
        weight_mem[16'h0E2D] <= 0;
        weight_mem[16'h0E2E] <= 0;
        weight_mem[16'h0E2F] <= 0;
        weight_mem[16'h0E30] <= 0;
        weight_mem[16'h0E31] <= 0;
        weight_mem[16'h0E32] <= 0;
        weight_mem[16'h0E33] <= 0;
        weight_mem[16'h0E34] <= 0;
        weight_mem[16'h0E35] <= 0;
        weight_mem[16'h0E36] <= 0;
        weight_mem[16'h0E37] <= 0;
        weight_mem[16'h0E38] <= 0;
        weight_mem[16'h0E39] <= 0;
        weight_mem[16'h0E3A] <= 0;
        weight_mem[16'h0E3B] <= 0;
        weight_mem[16'h0E3C] <= 0;
        weight_mem[16'h0E3D] <= 0;
        weight_mem[16'h0E3E] <= 0;
        weight_mem[16'h0E3F] <= 0;
        weight_mem[16'h0E40] <= 0;
        weight_mem[16'h0E41] <= 0;
        weight_mem[16'h0E42] <= 0;
        weight_mem[16'h0E43] <= 0;
        weight_mem[16'h0E44] <= 0;
        weight_mem[16'h0E45] <= 0;
        weight_mem[16'h0E46] <= 0;
        weight_mem[16'h0E47] <= 0;
        weight_mem[16'h0E48] <= 0;
        weight_mem[16'h0E49] <= 0;
        weight_mem[16'h0E4A] <= 0;
        weight_mem[16'h0E4B] <= 0;
        weight_mem[16'h0E4C] <= 0;
        weight_mem[16'h0E4D] <= 0;
        weight_mem[16'h0E4E] <= 0;
        weight_mem[16'h0E4F] <= 0;
        weight_mem[16'h0E50] <= 0;
        weight_mem[16'h0E51] <= 0;
        weight_mem[16'h0E52] <= 0;
        weight_mem[16'h0E53] <= 0;
        weight_mem[16'h0E54] <= 0;
        weight_mem[16'h0E55] <= 0;
        weight_mem[16'h0E56] <= 0;
        weight_mem[16'h0E57] <= 0;
        weight_mem[16'h0E58] <= 0;
        weight_mem[16'h0E59] <= 0;
        weight_mem[16'h0E5A] <= 0;
        weight_mem[16'h0E5B] <= 0;
        weight_mem[16'h0E5C] <= 0;
        weight_mem[16'h0E5D] <= 0;
        weight_mem[16'h0E5E] <= 0;
        weight_mem[16'h0E5F] <= 0;
        weight_mem[16'h0E60] <= 0;
        weight_mem[16'h0E61] <= 0;
        weight_mem[16'h0E62] <= 0;
        weight_mem[16'h0E63] <= 0;
        weight_mem[16'h0E64] <= 0;
        weight_mem[16'h0E65] <= 0;
        weight_mem[16'h0E66] <= 0;
        weight_mem[16'h0E67] <= 0;
        weight_mem[16'h0E68] <= 0;
        weight_mem[16'h0E69] <= 0;
        weight_mem[16'h0E6A] <= 0;
        weight_mem[16'h0E6B] <= 0;
        weight_mem[16'h0E6C] <= 0;
        weight_mem[16'h0E6D] <= 0;
        weight_mem[16'h0E6E] <= 0;
        weight_mem[16'h0E6F] <= 0;
        weight_mem[16'h0E70] <= 0;
        weight_mem[16'h0E71] <= 0;
        weight_mem[16'h0E72] <= 0;
        weight_mem[16'h0E73] <= 0;
        weight_mem[16'h0E74] <= 0;
        weight_mem[16'h0E75] <= 0;
        weight_mem[16'h0E76] <= 0;
        weight_mem[16'h0E77] <= 0;
        weight_mem[16'h0E78] <= 0;
        weight_mem[16'h0E79] <= 0;
        weight_mem[16'h0E7A] <= 0;
        weight_mem[16'h0E7B] <= 0;
        weight_mem[16'h0E7C] <= 0;
        weight_mem[16'h0E7D] <= 0;
        weight_mem[16'h0E7E] <= 0;
        weight_mem[16'h0E7F] <= 0;
        weight_mem[16'h0E80] <= 0;
        weight_mem[16'h0E81] <= 0;
        weight_mem[16'h0E82] <= 0;
        weight_mem[16'h0E83] <= 0;
        weight_mem[16'h0E84] <= 0;
        weight_mem[16'h0E85] <= 0;
        weight_mem[16'h0E86] <= 0;
        weight_mem[16'h0E87] <= 0;
        weight_mem[16'h0E88] <= 0;
        weight_mem[16'h0E89] <= 0;
        weight_mem[16'h0E8A] <= 0;
        weight_mem[16'h0E8B] <= 0;
        weight_mem[16'h0E8C] <= 0;
        weight_mem[16'h0E8D] <= 0;
        weight_mem[16'h0E8E] <= 0;
        weight_mem[16'h0E8F] <= 0;
        weight_mem[16'h0E90] <= 0;
        weight_mem[16'h0E91] <= 0;
        weight_mem[16'h0E92] <= 0;
        weight_mem[16'h0E93] <= 0;
        weight_mem[16'h0E94] <= 0;
        weight_mem[16'h0E95] <= 0;
        weight_mem[16'h0E96] <= 0;
        weight_mem[16'h0E97] <= 0;
        weight_mem[16'h0E98] <= 0;
        weight_mem[16'h0E99] <= 0;
        weight_mem[16'h0E9A] <= 0;
        weight_mem[16'h0E9B] <= 0;
        weight_mem[16'h0E9C] <= 0;
        weight_mem[16'h0E9D] <= 0;
        weight_mem[16'h0E9E] <= 0;
        weight_mem[16'h0E9F] <= 0;
        weight_mem[16'h0EA0] <= 0;
        weight_mem[16'h0EA1] <= 0;
        weight_mem[16'h0EA2] <= 0;
        weight_mem[16'h0EA3] <= 0;
        weight_mem[16'h0EA4] <= 0;
        weight_mem[16'h0EA5] <= 0;
        weight_mem[16'h0EA6] <= 0;
        weight_mem[16'h0EA7] <= 0;
        weight_mem[16'h0EA8] <= 0;
        weight_mem[16'h0EA9] <= 0;
        weight_mem[16'h0EAA] <= 0;
        weight_mem[16'h0EAB] <= 0;
        weight_mem[16'h0EAC] <= 0;
        weight_mem[16'h0EAD] <= 0;
        weight_mem[16'h0EAE] <= 0;
        weight_mem[16'h0EAF] <= 0;
        weight_mem[16'h0EB0] <= 0;
        weight_mem[16'h0EB1] <= 0;
        weight_mem[16'h0EB2] <= 0;
        weight_mem[16'h0EB3] <= 0;
        weight_mem[16'h0EB4] <= 0;
        weight_mem[16'h0EB5] <= 0;
        weight_mem[16'h0EB6] <= 0;
        weight_mem[16'h0EB7] <= 0;
        weight_mem[16'h0EB8] <= 0;
        weight_mem[16'h0EB9] <= 0;
        weight_mem[16'h0EBA] <= 0;
        weight_mem[16'h0EBB] <= 0;
        weight_mem[16'h0EBC] <= 0;
        weight_mem[16'h0EBD] <= 0;
        weight_mem[16'h0EBE] <= 0;
        weight_mem[16'h0EBF] <= 0;
        weight_mem[16'h0EC0] <= 0;
        weight_mem[16'h0EC1] <= 0;
        weight_mem[16'h0EC2] <= 0;
        weight_mem[16'h0EC3] <= 0;
        weight_mem[16'h0EC4] <= 0;
        weight_mem[16'h0EC5] <= 0;
        weight_mem[16'h0EC6] <= 0;
        weight_mem[16'h0EC7] <= 0;
        weight_mem[16'h0EC8] <= 0;
        weight_mem[16'h0EC9] <= 0;
        weight_mem[16'h0ECA] <= 0;
        weight_mem[16'h0ECB] <= 0;
        weight_mem[16'h0ECC] <= 0;
        weight_mem[16'h0ECD] <= 0;
        weight_mem[16'h0ECE] <= 0;
        weight_mem[16'h0ECF] <= 0;
        weight_mem[16'h0ED0] <= 0;
        weight_mem[16'h0ED1] <= 0;
        weight_mem[16'h0ED2] <= 0;
        weight_mem[16'h0ED3] <= 0;
        weight_mem[16'h0ED4] <= 0;
        weight_mem[16'h0ED5] <= 0;
        weight_mem[16'h0ED6] <= 0;
        weight_mem[16'h0ED7] <= 0;
        weight_mem[16'h0ED8] <= 0;
        weight_mem[16'h0ED9] <= 0;
        weight_mem[16'h0EDA] <= 0;
        weight_mem[16'h0EDB] <= 0;
        weight_mem[16'h0EDC] <= 0;
        weight_mem[16'h0EDD] <= 0;
        weight_mem[16'h0EDE] <= 0;
        weight_mem[16'h0EDF] <= 0;
        weight_mem[16'h0EE0] <= 0;
        weight_mem[16'h0EE1] <= 0;
        weight_mem[16'h0EE2] <= 0;
        weight_mem[16'h0EE3] <= 0;
        weight_mem[16'h0EE4] <= 0;
        weight_mem[16'h0EE5] <= 0;
        weight_mem[16'h0EE6] <= 0;
        weight_mem[16'h0EE7] <= 0;
        weight_mem[16'h0EE8] <= 0;
        weight_mem[16'h0EE9] <= 0;
        weight_mem[16'h0EEA] <= 0;
        weight_mem[16'h0EEB] <= 0;
        weight_mem[16'h0EEC] <= 0;
        weight_mem[16'h0EED] <= 0;
        weight_mem[16'h0EEE] <= 0;
        weight_mem[16'h0EEF] <= 0;
        weight_mem[16'h0EF0] <= 0;
        weight_mem[16'h0EF1] <= 0;
        weight_mem[16'h0EF2] <= 0;
        weight_mem[16'h0EF3] <= 0;
        weight_mem[16'h0EF4] <= 0;
        weight_mem[16'h0EF5] <= 0;
        weight_mem[16'h0EF6] <= 0;
        weight_mem[16'h0EF7] <= 0;
        weight_mem[16'h0EF8] <= 0;
        weight_mem[16'h0EF9] <= 0;
        weight_mem[16'h0EFA] <= 0;
        weight_mem[16'h0EFB] <= 0;
        weight_mem[16'h0EFC] <= 0;
        weight_mem[16'h0EFD] <= 0;
        weight_mem[16'h0EFE] <= 0;
        weight_mem[16'h0EFF] <= 0;
        weight_mem[16'h0F00] <= 0;
        weight_mem[16'h0F01] <= 0;
        weight_mem[16'h0F02] <= 0;
        weight_mem[16'h0F03] <= 0;
        weight_mem[16'h0F04] <= 0;
        weight_mem[16'h0F05] <= 0;
        weight_mem[16'h0F06] <= 0;
        weight_mem[16'h0F07] <= 0;
        weight_mem[16'h0F08] <= 0;
        weight_mem[16'h0F09] <= 0;
        weight_mem[16'h0F0A] <= 0;
        weight_mem[16'h0F0B] <= 0;
        weight_mem[16'h0F0C] <= 0;
        weight_mem[16'h0F0D] <= 0;
        weight_mem[16'h0F0E] <= 0;
        weight_mem[16'h0F0F] <= 0;
        weight_mem[16'h0F10] <= 0;
        weight_mem[16'h0F11] <= 0;
        weight_mem[16'h0F12] <= 0;
        weight_mem[16'h0F13] <= 0;
        weight_mem[16'h0F14] <= 0;
        weight_mem[16'h0F15] <= 0;
        weight_mem[16'h0F16] <= 0;
        weight_mem[16'h0F17] <= 0;
        weight_mem[16'h0F18] <= 0;
        weight_mem[16'h0F19] <= 0;
        weight_mem[16'h0F1A] <= 0;
        weight_mem[16'h0F1B] <= 0;
        weight_mem[16'h0F1C] <= 0;
        weight_mem[16'h0F1D] <= 0;
        weight_mem[16'h0F1E] <= 0;
        weight_mem[16'h0F1F] <= 0;
        weight_mem[16'h0F20] <= 0;
        weight_mem[16'h0F21] <= 0;
        weight_mem[16'h0F22] <= 0;
        weight_mem[16'h0F23] <= 0;
        weight_mem[16'h0F24] <= 0;
        weight_mem[16'h0F25] <= 0;
        weight_mem[16'h0F26] <= 0;
        weight_mem[16'h0F27] <= 0;
        weight_mem[16'h0F28] <= 0;
        weight_mem[16'h0F29] <= 0;
        weight_mem[16'h0F2A] <= 0;
        weight_mem[16'h0F2B] <= 0;
        weight_mem[16'h0F2C] <= 0;
        weight_mem[16'h0F2D] <= 0;
        weight_mem[16'h0F2E] <= 0;
        weight_mem[16'h0F2F] <= 0;
        weight_mem[16'h0F30] <= 0;
        weight_mem[16'h0F31] <= 0;
        weight_mem[16'h0F32] <= 0;
        weight_mem[16'h0F33] <= 0;
        weight_mem[16'h0F34] <= 0;
        weight_mem[16'h0F35] <= 0;
        weight_mem[16'h0F36] <= 0;
        weight_mem[16'h0F37] <= 0;
        weight_mem[16'h0F38] <= 0;
        weight_mem[16'h0F39] <= 0;
        weight_mem[16'h0F3A] <= 0;
        weight_mem[16'h0F3B] <= 0;
        weight_mem[16'h0F3C] <= 0;
        weight_mem[16'h0F3D] <= 0;
        weight_mem[16'h0F3E] <= 0;
        weight_mem[16'h0F3F] <= 0;
        weight_mem[16'h0F40] <= 0;
        weight_mem[16'h0F41] <= 0;
        weight_mem[16'h0F42] <= 0;
        weight_mem[16'h0F43] <= 0;
        weight_mem[16'h0F44] <= 0;
        weight_mem[16'h0F45] <= 0;
        weight_mem[16'h0F46] <= 0;
        weight_mem[16'h0F47] <= 0;
        weight_mem[16'h0F48] <= 0;
        weight_mem[16'h0F49] <= 0;
        weight_mem[16'h0F4A] <= 0;
        weight_mem[16'h0F4B] <= 0;
        weight_mem[16'h0F4C] <= 0;
        weight_mem[16'h0F4D] <= 0;
        weight_mem[16'h0F4E] <= 0;
        weight_mem[16'h0F4F] <= 0;
        weight_mem[16'h0F50] <= 0;
        weight_mem[16'h0F51] <= 0;
        weight_mem[16'h0F52] <= 0;
        weight_mem[16'h0F53] <= 0;
        weight_mem[16'h0F54] <= 0;
        weight_mem[16'h0F55] <= 0;
        weight_mem[16'h0F56] <= 0;
        weight_mem[16'h0F57] <= 0;
        weight_mem[16'h0F58] <= 0;
        weight_mem[16'h0F59] <= 0;
        weight_mem[16'h0F5A] <= 0;
        weight_mem[16'h0F5B] <= 0;
        weight_mem[16'h0F5C] <= 0;
        weight_mem[16'h0F5D] <= 0;
        weight_mem[16'h0F5E] <= 0;
        weight_mem[16'h0F5F] <= 0;
        weight_mem[16'h0F60] <= 0;
        weight_mem[16'h0F61] <= 0;
        weight_mem[16'h0F62] <= 0;
        weight_mem[16'h0F63] <= 0;
        weight_mem[16'h0F64] <= 0;
        weight_mem[16'h0F65] <= 0;
        weight_mem[16'h0F66] <= 0;
        weight_mem[16'h0F67] <= 0;
        weight_mem[16'h0F68] <= 0;
        weight_mem[16'h0F69] <= 0;
        weight_mem[16'h0F6A] <= 0;
        weight_mem[16'h0F6B] <= 0;
        weight_mem[16'h0F6C] <= 0;
        weight_mem[16'h0F6D] <= 0;
        weight_mem[16'h0F6E] <= 0;
        weight_mem[16'h0F6F] <= 0;
        weight_mem[16'h0F70] <= 0;
        weight_mem[16'h0F71] <= 0;
        weight_mem[16'h0F72] <= 0;
        weight_mem[16'h0F73] <= 0;
        weight_mem[16'h0F74] <= 0;
        weight_mem[16'h0F75] <= 0;
        weight_mem[16'h0F76] <= 0;
        weight_mem[16'h0F77] <= 0;
        weight_mem[16'h0F78] <= 0;
        weight_mem[16'h0F79] <= 0;
        weight_mem[16'h0F7A] <= 0;
        weight_mem[16'h0F7B] <= 0;
        weight_mem[16'h0F7C] <= 0;
        weight_mem[16'h0F7D] <= 0;
        weight_mem[16'h0F7E] <= 0;
        weight_mem[16'h0F7F] <= 0;
        weight_mem[16'h0F80] <= 0;
        weight_mem[16'h0F81] <= 0;
        weight_mem[16'h0F82] <= 0;
        weight_mem[16'h0F83] <= 0;
        weight_mem[16'h0F84] <= 0;
        weight_mem[16'h0F85] <= 0;
        weight_mem[16'h0F86] <= 0;
        weight_mem[16'h0F87] <= 0;
        weight_mem[16'h0F88] <= 0;
        weight_mem[16'h0F89] <= 0;
        weight_mem[16'h0F8A] <= 0;
        weight_mem[16'h0F8B] <= 0;
        weight_mem[16'h0F8C] <= 0;
        weight_mem[16'h0F8D] <= 0;
        weight_mem[16'h0F8E] <= 0;
        weight_mem[16'h0F8F] <= 0;
        weight_mem[16'h0F90] <= 0;
        weight_mem[16'h0F91] <= 0;
        weight_mem[16'h0F92] <= 0;
        weight_mem[16'h0F93] <= 0;
        weight_mem[16'h0F94] <= 0;
        weight_mem[16'h0F95] <= 0;
        weight_mem[16'h0F96] <= 0;
        weight_mem[16'h0F97] <= 0;
        weight_mem[16'h0F98] <= 0;
        weight_mem[16'h0F99] <= 0;
        weight_mem[16'h0F9A] <= 0;
        weight_mem[16'h0F9B] <= 0;
        weight_mem[16'h0F9C] <= 0;
        weight_mem[16'h0F9D] <= 0;
        weight_mem[16'h0F9E] <= 0;
        weight_mem[16'h0F9F] <= 0;
        weight_mem[16'h0FA0] <= 0;
        weight_mem[16'h0FA1] <= 0;
        weight_mem[16'h0FA2] <= 0;
        weight_mem[16'h0FA3] <= 0;
        weight_mem[16'h0FA4] <= 0;
        weight_mem[16'h0FA5] <= 0;
        weight_mem[16'h0FA6] <= 0;
        weight_mem[16'h0FA7] <= 0;
        weight_mem[16'h0FA8] <= 0;
        weight_mem[16'h0FA9] <= 0;
        weight_mem[16'h0FAA] <= 0;
        weight_mem[16'h0FAB] <= 0;
        weight_mem[16'h0FAC] <= 0;
        weight_mem[16'h0FAD] <= 0;
        weight_mem[16'h0FAE] <= 0;
        weight_mem[16'h0FAF] <= 0;

        // layer 1 neuron 8
        weight_mem[16'h1000] <= 0;
        weight_mem[16'h1001] <= 0;
        weight_mem[16'h1002] <= 0;
        weight_mem[16'h1003] <= 0;
        weight_mem[16'h1004] <= 0;
        weight_mem[16'h1005] <= 0;
        weight_mem[16'h1006] <= 0;
        weight_mem[16'h1007] <= 0;
        weight_mem[16'h1008] <= 0;
        weight_mem[16'h1009] <= 0;
        weight_mem[16'h100A] <= 0;
        weight_mem[16'h100B] <= 0;
        weight_mem[16'h100C] <= 0;
        weight_mem[16'h100D] <= 0;
        weight_mem[16'h100E] <= 0;
        weight_mem[16'h100F] <= 0;
        weight_mem[16'h1010] <= 0;
        weight_mem[16'h1011] <= 0;
        weight_mem[16'h1012] <= 0;
        weight_mem[16'h1013] <= 0;
        weight_mem[16'h1014] <= 0;
        weight_mem[16'h1015] <= 0;
        weight_mem[16'h1016] <= 0;
        weight_mem[16'h1017] <= 0;
        weight_mem[16'h1018] <= 0;
        weight_mem[16'h1019] <= 0;
        weight_mem[16'h101A] <= 0;
        weight_mem[16'h101B] <= 0;
        weight_mem[16'h101C] <= 0;
        weight_mem[16'h101D] <= 0;
        weight_mem[16'h101E] <= 0;
        weight_mem[16'h101F] <= 0;
        weight_mem[16'h1020] <= 0;
        weight_mem[16'h1021] <= 0;
        weight_mem[16'h1022] <= 0;
        weight_mem[16'h1023] <= 0;
        weight_mem[16'h1024] <= 0;
        weight_mem[16'h1025] <= 0;
        weight_mem[16'h1026] <= 0;
        weight_mem[16'h1027] <= 0;
        weight_mem[16'h1028] <= 0;
        weight_mem[16'h1029] <= 0;
        weight_mem[16'h102A] <= 0;
        weight_mem[16'h102B] <= 0;
        weight_mem[16'h102C] <= 0;
        weight_mem[16'h102D] <= 0;
        weight_mem[16'h102E] <= 0;
        weight_mem[16'h102F] <= 0;
        weight_mem[16'h1030] <= 0;
        weight_mem[16'h1031] <= 0;
        weight_mem[16'h1032] <= 0;
        weight_mem[16'h1033] <= 0;
        weight_mem[16'h1034] <= 0;
        weight_mem[16'h1035] <= 0;
        weight_mem[16'h1036] <= 0;
        weight_mem[16'h1037] <= 0;
        weight_mem[16'h1038] <= 0;
        weight_mem[16'h1039] <= 0;
        weight_mem[16'h103A] <= 0;
        weight_mem[16'h103B] <= 0;
        weight_mem[16'h103C] <= 0;
        weight_mem[16'h103D] <= 0;
        weight_mem[16'h103E] <= 0;
        weight_mem[16'h103F] <= 0;
        weight_mem[16'h1040] <= 0;
        weight_mem[16'h1041] <= 0;
        weight_mem[16'h1042] <= 0;
        weight_mem[16'h1043] <= 0;
        weight_mem[16'h1044] <= 0;
        weight_mem[16'h1045] <= 0;
        weight_mem[16'h1046] <= 0;
        weight_mem[16'h1047] <= 0;
        weight_mem[16'h1048] <= 0;
        weight_mem[16'h1049] <= 0;
        weight_mem[16'h104A] <= 0;
        weight_mem[16'h104B] <= 0;
        weight_mem[16'h104C] <= 0;
        weight_mem[16'h104D] <= 0;
        weight_mem[16'h104E] <= 0;
        weight_mem[16'h104F] <= 0;
        weight_mem[16'h1050] <= 0;
        weight_mem[16'h1051] <= 0;
        weight_mem[16'h1052] <= 0;
        weight_mem[16'h1053] <= 0;
        weight_mem[16'h1054] <= 0;
        weight_mem[16'h1055] <= 0;
        weight_mem[16'h1056] <= 0;
        weight_mem[16'h1057] <= 0;
        weight_mem[16'h1058] <= 0;
        weight_mem[16'h1059] <= 0;
        weight_mem[16'h105A] <= 0;
        weight_mem[16'h105B] <= 0;
        weight_mem[16'h105C] <= 0;
        weight_mem[16'h105D] <= 0;
        weight_mem[16'h105E] <= 0;
        weight_mem[16'h105F] <= 0;
        weight_mem[16'h1060] <= 0;
        weight_mem[16'h1061] <= 0;
        weight_mem[16'h1062] <= 0;
        weight_mem[16'h1063] <= 0;
        weight_mem[16'h1064] <= 0;
        weight_mem[16'h1065] <= 0;
        weight_mem[16'h1066] <= 0;
        weight_mem[16'h1067] <= 0;
        weight_mem[16'h1068] <= 0;
        weight_mem[16'h1069] <= 0;
        weight_mem[16'h106A] <= 0;
        weight_mem[16'h106B] <= 0;
        weight_mem[16'h106C] <= 0;
        weight_mem[16'h106D] <= 0;
        weight_mem[16'h106E] <= 0;
        weight_mem[16'h106F] <= 0;
        weight_mem[16'h1070] <= 0;
        weight_mem[16'h1071] <= 0;
        weight_mem[16'h1072] <= 0;
        weight_mem[16'h1073] <= 0;
        weight_mem[16'h1074] <= 0;
        weight_mem[16'h1075] <= 0;
        weight_mem[16'h1076] <= 0;
        weight_mem[16'h1077] <= 0;
        weight_mem[16'h1078] <= 0;
        weight_mem[16'h1079] <= 0;
        weight_mem[16'h107A] <= 0;
        weight_mem[16'h107B] <= 0;
        weight_mem[16'h107C] <= 0;
        weight_mem[16'h107D] <= 0;
        weight_mem[16'h107E] <= 0;
        weight_mem[16'h107F] <= 0;
        weight_mem[16'h1080] <= 0;
        weight_mem[16'h1081] <= 0;
        weight_mem[16'h1082] <= 0;
        weight_mem[16'h1083] <= 0;
        weight_mem[16'h1084] <= 0;
        weight_mem[16'h1085] <= 0;
        weight_mem[16'h1086] <= 0;
        weight_mem[16'h1087] <= 0;
        weight_mem[16'h1088] <= 0;
        weight_mem[16'h1089] <= 0;
        weight_mem[16'h108A] <= 0;
        weight_mem[16'h108B] <= 0;
        weight_mem[16'h108C] <= 0;
        weight_mem[16'h108D] <= 0;
        weight_mem[16'h108E] <= 0;
        weight_mem[16'h108F] <= 0;
        weight_mem[16'h1090] <= 0;
        weight_mem[16'h1091] <= 0;
        weight_mem[16'h1092] <= 0;
        weight_mem[16'h1093] <= 0;
        weight_mem[16'h1094] <= 0;
        weight_mem[16'h1095] <= 0;
        weight_mem[16'h1096] <= 0;
        weight_mem[16'h1097] <= 0;
        weight_mem[16'h1098] <= 0;
        weight_mem[16'h1099] <= 0;
        weight_mem[16'h109A] <= 0;
        weight_mem[16'h109B] <= 0;
        weight_mem[16'h109C] <= 0;
        weight_mem[16'h109D] <= 0;
        weight_mem[16'h109E] <= 0;
        weight_mem[16'h109F] <= 0;
        weight_mem[16'h10A0] <= 0;
        weight_mem[16'h10A1] <= 0;
        weight_mem[16'h10A2] <= 0;
        weight_mem[16'h10A3] <= 0;
        weight_mem[16'h10A4] <= 0;
        weight_mem[16'h10A5] <= 0;
        weight_mem[16'h10A6] <= 0;
        weight_mem[16'h10A7] <= 0;
        weight_mem[16'h10A8] <= 0;
        weight_mem[16'h10A9] <= 0;
        weight_mem[16'h10AA] <= 0;
        weight_mem[16'h10AB] <= 0;
        weight_mem[16'h10AC] <= 0;
        weight_mem[16'h10AD] <= 0;
        weight_mem[16'h10AE] <= 0;
        weight_mem[16'h10AF] <= 0;
        weight_mem[16'h10B0] <= 0;
        weight_mem[16'h10B1] <= 0;
        weight_mem[16'h10B2] <= 0;
        weight_mem[16'h10B3] <= 0;
        weight_mem[16'h10B4] <= 0;
        weight_mem[16'h10B5] <= 0;
        weight_mem[16'h10B6] <= 0;
        weight_mem[16'h10B7] <= 0;
        weight_mem[16'h10B8] <= 0;
        weight_mem[16'h10B9] <= 0;
        weight_mem[16'h10BA] <= 0;
        weight_mem[16'h10BB] <= 0;
        weight_mem[16'h10BC] <= 0;
        weight_mem[16'h10BD] <= 0;
        weight_mem[16'h10BE] <= 0;
        weight_mem[16'h10BF] <= 0;
        weight_mem[16'h10C0] <= 0;
        weight_mem[16'h10C1] <= 0;
        weight_mem[16'h10C2] <= 0;
        weight_mem[16'h10C3] <= 0;
        weight_mem[16'h10C4] <= 0;
        weight_mem[16'h10C5] <= 0;
        weight_mem[16'h10C6] <= 0;
        weight_mem[16'h10C7] <= 0;
        weight_mem[16'h10C8] <= 0;
        weight_mem[16'h10C9] <= 0;
        weight_mem[16'h10CA] <= 0;
        weight_mem[16'h10CB] <= 0;
        weight_mem[16'h10CC] <= 0;
        weight_mem[16'h10CD] <= 0;
        weight_mem[16'h10CE] <= 0;
        weight_mem[16'h10CF] <= 0;
        weight_mem[16'h10D0] <= 0;
        weight_mem[16'h10D1] <= 0;
        weight_mem[16'h10D2] <= 0;
        weight_mem[16'h10D3] <= 0;
        weight_mem[16'h10D4] <= 0;
        weight_mem[16'h10D5] <= 0;
        weight_mem[16'h10D6] <= 0;
        weight_mem[16'h10D7] <= 0;
        weight_mem[16'h10D8] <= 0;
        weight_mem[16'h10D9] <= 0;
        weight_mem[16'h10DA] <= 0;
        weight_mem[16'h10DB] <= 0;
        weight_mem[16'h10DC] <= 0;
        weight_mem[16'h10DD] <= 0;
        weight_mem[16'h10DE] <= 0;
        weight_mem[16'h10DF] <= 0;
        weight_mem[16'h10E0] <= 0;
        weight_mem[16'h10E1] <= 0;
        weight_mem[16'h10E2] <= 0;
        weight_mem[16'h10E3] <= 0;
        weight_mem[16'h10E4] <= 0;
        weight_mem[16'h10E5] <= 0;
        weight_mem[16'h10E6] <= 0;
        weight_mem[16'h10E7] <= 0;
        weight_mem[16'h10E8] <= 0;
        weight_mem[16'h10E9] <= 0;
        weight_mem[16'h10EA] <= 0;
        weight_mem[16'h10EB] <= 0;
        weight_mem[16'h10EC] <= 0;
        weight_mem[16'h10ED] <= 0;
        weight_mem[16'h10EE] <= 0;
        weight_mem[16'h10EF] <= 0;
        weight_mem[16'h10F0] <= 0;
        weight_mem[16'h10F1] <= 0;
        weight_mem[16'h10F2] <= 0;
        weight_mem[16'h10F3] <= 0;
        weight_mem[16'h10F4] <= 0;
        weight_mem[16'h10F5] <= 0;
        weight_mem[16'h10F6] <= 0;
        weight_mem[16'h10F7] <= 0;
        weight_mem[16'h10F8] <= 0;
        weight_mem[16'h10F9] <= 0;
        weight_mem[16'h10FA] <= 0;
        weight_mem[16'h10FB] <= 0;
        weight_mem[16'h10FC] <= 0;
        weight_mem[16'h10FD] <= 0;
        weight_mem[16'h10FE] <= 0;
        weight_mem[16'h10FF] <= 0;
        weight_mem[16'h1100] <= 0;
        weight_mem[16'h1101] <= 0;
        weight_mem[16'h1102] <= 0;
        weight_mem[16'h1103] <= 0;
        weight_mem[16'h1104] <= 0;
        weight_mem[16'h1105] <= 0;
        weight_mem[16'h1106] <= 0;
        weight_mem[16'h1107] <= 0;
        weight_mem[16'h1108] <= 0;
        weight_mem[16'h1109] <= 0;
        weight_mem[16'h110A] <= 0;
        weight_mem[16'h110B] <= 0;
        weight_mem[16'h110C] <= 0;
        weight_mem[16'h110D] <= 0;
        weight_mem[16'h110E] <= 0;
        weight_mem[16'h110F] <= 0;
        weight_mem[16'h1110] <= 0;
        weight_mem[16'h1111] <= 0;
        weight_mem[16'h1112] <= 0;
        weight_mem[16'h1113] <= 0;
        weight_mem[16'h1114] <= 0;
        weight_mem[16'h1115] <= 0;
        weight_mem[16'h1116] <= 0;
        weight_mem[16'h1117] <= 0;
        weight_mem[16'h1118] <= 0;
        weight_mem[16'h1119] <= 0;
        weight_mem[16'h111A] <= 0;
        weight_mem[16'h111B] <= 0;
        weight_mem[16'h111C] <= 0;
        weight_mem[16'h111D] <= 0;
        weight_mem[16'h111E] <= 0;
        weight_mem[16'h111F] <= 0;
        weight_mem[16'h1120] <= 0;
        weight_mem[16'h1121] <= 0;
        weight_mem[16'h1122] <= 0;
        weight_mem[16'h1123] <= 0;
        weight_mem[16'h1124] <= 0;
        weight_mem[16'h1125] <= 0;
        weight_mem[16'h1126] <= 0;
        weight_mem[16'h1127] <= 0;
        weight_mem[16'h1128] <= 0;
        weight_mem[16'h1129] <= 0;
        weight_mem[16'h112A] <= 0;
        weight_mem[16'h112B] <= 0;
        weight_mem[16'h112C] <= 0;
        weight_mem[16'h112D] <= 0;
        weight_mem[16'h112E] <= 0;
        weight_mem[16'h112F] <= 0;
        weight_mem[16'h1130] <= 0;
        weight_mem[16'h1131] <= 0;
        weight_mem[16'h1132] <= 0;
        weight_mem[16'h1133] <= 0;
        weight_mem[16'h1134] <= 0;
        weight_mem[16'h1135] <= 0;
        weight_mem[16'h1136] <= 0;
        weight_mem[16'h1137] <= 0;
        weight_mem[16'h1138] <= 0;
        weight_mem[16'h1139] <= 0;
        weight_mem[16'h113A] <= 0;
        weight_mem[16'h113B] <= 0;
        weight_mem[16'h113C] <= 0;
        weight_mem[16'h113D] <= 0;
        weight_mem[16'h113E] <= 0;
        weight_mem[16'h113F] <= 0;
        weight_mem[16'h1140] <= 0;
        weight_mem[16'h1141] <= 0;
        weight_mem[16'h1142] <= 0;
        weight_mem[16'h1143] <= 0;
        weight_mem[16'h1144] <= 0;
        weight_mem[16'h1145] <= 0;
        weight_mem[16'h1146] <= 0;
        weight_mem[16'h1147] <= 0;
        weight_mem[16'h1148] <= 0;
        weight_mem[16'h1149] <= 0;
        weight_mem[16'h114A] <= 0;
        weight_mem[16'h114B] <= 0;
        weight_mem[16'h114C] <= 0;
        weight_mem[16'h114D] <= 0;
        weight_mem[16'h114E] <= 0;
        weight_mem[16'h114F] <= 0;
        weight_mem[16'h1150] <= 0;
        weight_mem[16'h1151] <= 0;
        weight_mem[16'h1152] <= 0;
        weight_mem[16'h1153] <= 0;
        weight_mem[16'h1154] <= 0;
        weight_mem[16'h1155] <= 0;
        weight_mem[16'h1156] <= 0;
        weight_mem[16'h1157] <= 0;
        weight_mem[16'h1158] <= 0;
        weight_mem[16'h1159] <= 0;
        weight_mem[16'h115A] <= 0;
        weight_mem[16'h115B] <= 0;
        weight_mem[16'h115C] <= 0;
        weight_mem[16'h115D] <= 0;
        weight_mem[16'h115E] <= 0;
        weight_mem[16'h115F] <= 0;
        weight_mem[16'h1160] <= 0;
        weight_mem[16'h1161] <= 0;
        weight_mem[16'h1162] <= 0;
        weight_mem[16'h1163] <= 0;
        weight_mem[16'h1164] <= 0;
        weight_mem[16'h1165] <= 0;
        weight_mem[16'h1166] <= 0;
        weight_mem[16'h1167] <= 0;
        weight_mem[16'h1168] <= 0;
        weight_mem[16'h1169] <= 0;
        weight_mem[16'h116A] <= 0;
        weight_mem[16'h116B] <= 0;
        weight_mem[16'h116C] <= 0;
        weight_mem[16'h116D] <= 0;
        weight_mem[16'h116E] <= 0;
        weight_mem[16'h116F] <= 0;
        weight_mem[16'h1170] <= 0;
        weight_mem[16'h1171] <= 0;
        weight_mem[16'h1172] <= 0;
        weight_mem[16'h1173] <= 0;
        weight_mem[16'h1174] <= 0;
        weight_mem[16'h1175] <= 0;
        weight_mem[16'h1176] <= 0;
        weight_mem[16'h1177] <= 0;
        weight_mem[16'h1178] <= 0;
        weight_mem[16'h1179] <= 0;
        weight_mem[16'h117A] <= 0;
        weight_mem[16'h117B] <= 0;
        weight_mem[16'h117C] <= 0;
        weight_mem[16'h117D] <= 0;
        weight_mem[16'h117E] <= 0;
        weight_mem[16'h117F] <= 0;
        weight_mem[16'h1180] <= 0;
        weight_mem[16'h1181] <= 0;
        weight_mem[16'h1182] <= 0;
        weight_mem[16'h1183] <= 0;
        weight_mem[16'h1184] <= 0;
        weight_mem[16'h1185] <= 0;
        weight_mem[16'h1186] <= 0;
        weight_mem[16'h1187] <= 0;
        weight_mem[16'h1188] <= 0;
        weight_mem[16'h1189] <= 0;
        weight_mem[16'h118A] <= 0;
        weight_mem[16'h118B] <= 0;
        weight_mem[16'h118C] <= 0;
        weight_mem[16'h118D] <= 0;
        weight_mem[16'h118E] <= 0;
        weight_mem[16'h118F] <= 0;
        weight_mem[16'h1190] <= 0;
        weight_mem[16'h1191] <= 0;
        weight_mem[16'h1192] <= 0;
        weight_mem[16'h1193] <= 0;
        weight_mem[16'h1194] <= 0;
        weight_mem[16'h1195] <= 0;
        weight_mem[16'h1196] <= 0;
        weight_mem[16'h1197] <= 0;
        weight_mem[16'h1198] <= 0;
        weight_mem[16'h1199] <= 0;
        weight_mem[16'h119A] <= 0;
        weight_mem[16'h119B] <= 0;
        weight_mem[16'h119C] <= 0;
        weight_mem[16'h119D] <= 0;
        weight_mem[16'h119E] <= 0;
        weight_mem[16'h119F] <= 0;
        weight_mem[16'h11A0] <= 0;
        weight_mem[16'h11A1] <= 0;
        weight_mem[16'h11A2] <= 0;
        weight_mem[16'h11A3] <= 0;
        weight_mem[16'h11A4] <= 0;
        weight_mem[16'h11A5] <= 0;
        weight_mem[16'h11A6] <= 0;
        weight_mem[16'h11A7] <= 0;
        weight_mem[16'h11A8] <= 0;
        weight_mem[16'h11A9] <= 0;
        weight_mem[16'h11AA] <= 0;
        weight_mem[16'h11AB] <= 0;
        weight_mem[16'h11AC] <= 0;
        weight_mem[16'h11AD] <= 0;
        weight_mem[16'h11AE] <= 0;
        weight_mem[16'h11AF] <= 0;

        // layer 1 neuron 9
        weight_mem[16'h1200] <= 0;
        weight_mem[16'h1201] <= 0;
        weight_mem[16'h1202] <= 0;
        weight_mem[16'h1203] <= 0;
        weight_mem[16'h1204] <= 0;
        weight_mem[16'h1205] <= 0;
        weight_mem[16'h1206] <= 0;
        weight_mem[16'h1207] <= 0;
        weight_mem[16'h1208] <= 0;
        weight_mem[16'h1209] <= 0;
        weight_mem[16'h120A] <= 0;
        weight_mem[16'h120B] <= 0;
        weight_mem[16'h120C] <= 0;
        weight_mem[16'h120D] <= 0;
        weight_mem[16'h120E] <= 0;
        weight_mem[16'h120F] <= 0;
        weight_mem[16'h1210] <= 0;
        weight_mem[16'h1211] <= 0;
        weight_mem[16'h1212] <= 0;
        weight_mem[16'h1213] <= 0;
        weight_mem[16'h1214] <= 0;
        weight_mem[16'h1215] <= 0;
        weight_mem[16'h1216] <= 0;
        weight_mem[16'h1217] <= 0;
        weight_mem[16'h1218] <= 0;
        weight_mem[16'h1219] <= 0;
        weight_mem[16'h121A] <= 0;
        weight_mem[16'h121B] <= 0;
        weight_mem[16'h121C] <= 0;
        weight_mem[16'h121D] <= 0;
        weight_mem[16'h121E] <= 0;
        weight_mem[16'h121F] <= 0;
        weight_mem[16'h1220] <= 0;
        weight_mem[16'h1221] <= 0;
        weight_mem[16'h1222] <= 0;
        weight_mem[16'h1223] <= 0;
        weight_mem[16'h1224] <= 0;
        weight_mem[16'h1225] <= 0;
        weight_mem[16'h1226] <= 0;
        weight_mem[16'h1227] <= 0;
        weight_mem[16'h1228] <= 0;
        weight_mem[16'h1229] <= 0;
        weight_mem[16'h122A] <= 0;
        weight_mem[16'h122B] <= 0;
        weight_mem[16'h122C] <= 0;
        weight_mem[16'h122D] <= 0;
        weight_mem[16'h122E] <= 0;
        weight_mem[16'h122F] <= 0;
        weight_mem[16'h1230] <= 0;
        weight_mem[16'h1231] <= 0;
        weight_mem[16'h1232] <= 0;
        weight_mem[16'h1233] <= 0;
        weight_mem[16'h1234] <= 0;
        weight_mem[16'h1235] <= 0;
        weight_mem[16'h1236] <= 0;
        weight_mem[16'h1237] <= 0;
        weight_mem[16'h1238] <= 0;
        weight_mem[16'h1239] <= 0;
        weight_mem[16'h123A] <= 0;
        weight_mem[16'h123B] <= 0;
        weight_mem[16'h123C] <= 0;
        weight_mem[16'h123D] <= 0;
        weight_mem[16'h123E] <= 0;
        weight_mem[16'h123F] <= 0;
        weight_mem[16'h1240] <= 0;
        weight_mem[16'h1241] <= 0;
        weight_mem[16'h1242] <= 0;
        weight_mem[16'h1243] <= 0;
        weight_mem[16'h1244] <= 0;
        weight_mem[16'h1245] <= 0;
        weight_mem[16'h1246] <= 0;
        weight_mem[16'h1247] <= 0;
        weight_mem[16'h1248] <= 0;
        weight_mem[16'h1249] <= 0;
        weight_mem[16'h124A] <= 0;
        weight_mem[16'h124B] <= 0;
        weight_mem[16'h124C] <= 0;
        weight_mem[16'h124D] <= 0;
        weight_mem[16'h124E] <= 0;
        weight_mem[16'h124F] <= 0;
        weight_mem[16'h1250] <= 0;
        weight_mem[16'h1251] <= 0;
        weight_mem[16'h1252] <= 0;
        weight_mem[16'h1253] <= 0;
        weight_mem[16'h1254] <= 0;
        weight_mem[16'h1255] <= 0;
        weight_mem[16'h1256] <= 0;
        weight_mem[16'h1257] <= 0;
        weight_mem[16'h1258] <= 0;
        weight_mem[16'h1259] <= 0;
        weight_mem[16'h125A] <= 0;
        weight_mem[16'h125B] <= 0;
        weight_mem[16'h125C] <= 0;
        weight_mem[16'h125D] <= 0;
        weight_mem[16'h125E] <= 0;
        weight_mem[16'h125F] <= 0;
        weight_mem[16'h1260] <= 0;
        weight_mem[16'h1261] <= 0;
        weight_mem[16'h1262] <= 0;
        weight_mem[16'h1263] <= 0;
        weight_mem[16'h1264] <= 0;
        weight_mem[16'h1265] <= 0;
        weight_mem[16'h1266] <= 0;
        weight_mem[16'h1267] <= 0;
        weight_mem[16'h1268] <= 0;
        weight_mem[16'h1269] <= 0;
        weight_mem[16'h126A] <= 0;
        weight_mem[16'h126B] <= 0;
        weight_mem[16'h126C] <= 0;
        weight_mem[16'h126D] <= 0;
        weight_mem[16'h126E] <= 0;
        weight_mem[16'h126F] <= 0;
        weight_mem[16'h1270] <= 0;
        weight_mem[16'h1271] <= 0;
        weight_mem[16'h1272] <= 0;
        weight_mem[16'h1273] <= 0;
        weight_mem[16'h1274] <= 0;
        weight_mem[16'h1275] <= 0;
        weight_mem[16'h1276] <= 0;
        weight_mem[16'h1277] <= 0;
        weight_mem[16'h1278] <= 0;
        weight_mem[16'h1279] <= 0;
        weight_mem[16'h127A] <= 0;
        weight_mem[16'h127B] <= 0;
        weight_mem[16'h127C] <= 0;
        weight_mem[16'h127D] <= 0;
        weight_mem[16'h127E] <= 0;
        weight_mem[16'h127F] <= 0;
        weight_mem[16'h1280] <= 0;
        weight_mem[16'h1281] <= 0;
        weight_mem[16'h1282] <= 0;
        weight_mem[16'h1283] <= 0;
        weight_mem[16'h1284] <= 0;
        weight_mem[16'h1285] <= 0;
        weight_mem[16'h1286] <= 0;
        weight_mem[16'h1287] <= 0;
        weight_mem[16'h1288] <= 0;
        weight_mem[16'h1289] <= 0;
        weight_mem[16'h128A] <= 0;
        weight_mem[16'h128B] <= 0;
        weight_mem[16'h128C] <= 0;
        weight_mem[16'h128D] <= 0;
        weight_mem[16'h128E] <= 0;
        weight_mem[16'h128F] <= 0;
        weight_mem[16'h1290] <= 0;
        weight_mem[16'h1291] <= 0;
        weight_mem[16'h1292] <= 0;
        weight_mem[16'h1293] <= 0;
        weight_mem[16'h1294] <= 0;
        weight_mem[16'h1295] <= 0;
        weight_mem[16'h1296] <= 0;
        weight_mem[16'h1297] <= 0;
        weight_mem[16'h1298] <= 0;
        weight_mem[16'h1299] <= 0;
        weight_mem[16'h129A] <= 0;
        weight_mem[16'h129B] <= 0;
        weight_mem[16'h129C] <= 0;
        weight_mem[16'h129D] <= 0;
        weight_mem[16'h129E] <= 0;
        weight_mem[16'h129F] <= 0;
        weight_mem[16'h12A0] <= 0;
        weight_mem[16'h12A1] <= 0;
        weight_mem[16'h12A2] <= 0;
        weight_mem[16'h12A3] <= 0;
        weight_mem[16'h12A4] <= 0;
        weight_mem[16'h12A5] <= 0;
        weight_mem[16'h12A6] <= 0;
        weight_mem[16'h12A7] <= 0;
        weight_mem[16'h12A8] <= 0;
        weight_mem[16'h12A9] <= 0;
        weight_mem[16'h12AA] <= 0;
        weight_mem[16'h12AB] <= 0;
        weight_mem[16'h12AC] <= 0;
        weight_mem[16'h12AD] <= 0;
        weight_mem[16'h12AE] <= 0;
        weight_mem[16'h12AF] <= 0;
        weight_mem[16'h12B0] <= 0;
        weight_mem[16'h12B1] <= 0;
        weight_mem[16'h12B2] <= 0;
        weight_mem[16'h12B3] <= 0;
        weight_mem[16'h12B4] <= 0;
        weight_mem[16'h12B5] <= 0;
        weight_mem[16'h12B6] <= 0;
        weight_mem[16'h12B7] <= 0;
        weight_mem[16'h12B8] <= 0;
        weight_mem[16'h12B9] <= 0;
        weight_mem[16'h12BA] <= 0;
        weight_mem[16'h12BB] <= 0;
        weight_mem[16'h12BC] <= 0;
        weight_mem[16'h12BD] <= 0;
        weight_mem[16'h12BE] <= 0;
        weight_mem[16'h12BF] <= 0;
        weight_mem[16'h12C0] <= 0;
        weight_mem[16'h12C1] <= 0;
        weight_mem[16'h12C2] <= 0;
        weight_mem[16'h12C3] <= 0;
        weight_mem[16'h12C4] <= 0;
        weight_mem[16'h12C5] <= 0;
        weight_mem[16'h12C6] <= 0;
        weight_mem[16'h12C7] <= 0;
        weight_mem[16'h12C8] <= 0;
        weight_mem[16'h12C9] <= 0;
        weight_mem[16'h12CA] <= 0;
        weight_mem[16'h12CB] <= 0;
        weight_mem[16'h12CC] <= 0;
        weight_mem[16'h12CD] <= 0;
        weight_mem[16'h12CE] <= 0;
        weight_mem[16'h12CF] <= 0;
        weight_mem[16'h12D0] <= 0;
        weight_mem[16'h12D1] <= 0;
        weight_mem[16'h12D2] <= 0;
        weight_mem[16'h12D3] <= 0;
        weight_mem[16'h12D4] <= 0;
        weight_mem[16'h12D5] <= 0;
        weight_mem[16'h12D6] <= 0;
        weight_mem[16'h12D7] <= 0;
        weight_mem[16'h12D8] <= 0;
        weight_mem[16'h12D9] <= 0;
        weight_mem[16'h12DA] <= 0;
        weight_mem[16'h12DB] <= 0;
        weight_mem[16'h12DC] <= 0;
        weight_mem[16'h12DD] <= 0;
        weight_mem[16'h12DE] <= 0;
        weight_mem[16'h12DF] <= 0;
        weight_mem[16'h12E0] <= 0;
        weight_mem[16'h12E1] <= 0;
        weight_mem[16'h12E2] <= 0;
        weight_mem[16'h12E3] <= 0;
        weight_mem[16'h12E4] <= 0;
        weight_mem[16'h12E5] <= 0;
        weight_mem[16'h12E6] <= 0;
        weight_mem[16'h12E7] <= 0;
        weight_mem[16'h12E8] <= 0;
        weight_mem[16'h12E9] <= 0;
        weight_mem[16'h12EA] <= 0;
        weight_mem[16'h12EB] <= 0;
        weight_mem[16'h12EC] <= 0;
        weight_mem[16'h12ED] <= 0;
        weight_mem[16'h12EE] <= 0;
        weight_mem[16'h12EF] <= 0;
        weight_mem[16'h12F0] <= 0;
        weight_mem[16'h12F1] <= 0;
        weight_mem[16'h12F2] <= 0;
        weight_mem[16'h12F3] <= 0;
        weight_mem[16'h12F4] <= 0;
        weight_mem[16'h12F5] <= 0;
        weight_mem[16'h12F6] <= 0;
        weight_mem[16'h12F7] <= 0;
        weight_mem[16'h12F8] <= 0;
        weight_mem[16'h12F9] <= 0;
        weight_mem[16'h12FA] <= 0;
        weight_mem[16'h12FB] <= 0;
        weight_mem[16'h12FC] <= 0;
        weight_mem[16'h12FD] <= 0;
        weight_mem[16'h12FE] <= 0;
        weight_mem[16'h12FF] <= 0;
        weight_mem[16'h1300] <= 0;
        weight_mem[16'h1301] <= 0;
        weight_mem[16'h1302] <= 0;
        weight_mem[16'h1303] <= 0;
        weight_mem[16'h1304] <= 0;
        weight_mem[16'h1305] <= 0;
        weight_mem[16'h1306] <= 0;
        weight_mem[16'h1307] <= 0;
        weight_mem[16'h1308] <= 0;
        weight_mem[16'h1309] <= 0;
        weight_mem[16'h130A] <= 0;
        weight_mem[16'h130B] <= 0;
        weight_mem[16'h130C] <= 0;
        weight_mem[16'h130D] <= 0;
        weight_mem[16'h130E] <= 0;
        weight_mem[16'h130F] <= 0;
        weight_mem[16'h1310] <= 0;
        weight_mem[16'h1311] <= 0;
        weight_mem[16'h1312] <= 0;
        weight_mem[16'h1313] <= 0;
        weight_mem[16'h1314] <= 0;
        weight_mem[16'h1315] <= 0;
        weight_mem[16'h1316] <= 0;
        weight_mem[16'h1317] <= 0;
        weight_mem[16'h1318] <= 0;
        weight_mem[16'h1319] <= 0;
        weight_mem[16'h131A] <= 0;
        weight_mem[16'h131B] <= 0;
        weight_mem[16'h131C] <= 0;
        weight_mem[16'h131D] <= 0;
        weight_mem[16'h131E] <= 0;
        weight_mem[16'h131F] <= 0;
        weight_mem[16'h1320] <= 0;
        weight_mem[16'h1321] <= 0;
        weight_mem[16'h1322] <= 0;
        weight_mem[16'h1323] <= 0;
        weight_mem[16'h1324] <= 0;
        weight_mem[16'h1325] <= 0;
        weight_mem[16'h1326] <= 0;
        weight_mem[16'h1327] <= 0;
        weight_mem[16'h1328] <= 0;
        weight_mem[16'h1329] <= 0;
        weight_mem[16'h132A] <= 0;
        weight_mem[16'h132B] <= 0;
        weight_mem[16'h132C] <= 0;
        weight_mem[16'h132D] <= 0;
        weight_mem[16'h132E] <= 0;
        weight_mem[16'h132F] <= 0;
        weight_mem[16'h1330] <= 0;
        weight_mem[16'h1331] <= 0;
        weight_mem[16'h1332] <= 0;
        weight_mem[16'h1333] <= 0;
        weight_mem[16'h1334] <= 0;
        weight_mem[16'h1335] <= 0;
        weight_mem[16'h1336] <= 0;
        weight_mem[16'h1337] <= 0;
        weight_mem[16'h1338] <= 0;
        weight_mem[16'h1339] <= 0;
        weight_mem[16'h133A] <= 0;
        weight_mem[16'h133B] <= 0;
        weight_mem[16'h133C] <= 0;
        weight_mem[16'h133D] <= 0;
        weight_mem[16'h133E] <= 0;
        weight_mem[16'h133F] <= 0;
        weight_mem[16'h1340] <= 0;
        weight_mem[16'h1341] <= 0;
        weight_mem[16'h1342] <= 0;
        weight_mem[16'h1343] <= 0;
        weight_mem[16'h1344] <= 0;
        weight_mem[16'h1345] <= 0;
        weight_mem[16'h1346] <= 0;
        weight_mem[16'h1347] <= 0;
        weight_mem[16'h1348] <= 0;
        weight_mem[16'h1349] <= 0;
        weight_mem[16'h134A] <= 0;
        weight_mem[16'h134B] <= 0;
        weight_mem[16'h134C] <= 0;
        weight_mem[16'h134D] <= 0;
        weight_mem[16'h134E] <= 0;
        weight_mem[16'h134F] <= 0;
        weight_mem[16'h1350] <= 0;
        weight_mem[16'h1351] <= 0;
        weight_mem[16'h1352] <= 0;
        weight_mem[16'h1353] <= 0;
        weight_mem[16'h1354] <= 0;
        weight_mem[16'h1355] <= 0;
        weight_mem[16'h1356] <= 0;
        weight_mem[16'h1357] <= 0;
        weight_mem[16'h1358] <= 0;
        weight_mem[16'h1359] <= 0;
        weight_mem[16'h135A] <= 0;
        weight_mem[16'h135B] <= 0;
        weight_mem[16'h135C] <= 0;
        weight_mem[16'h135D] <= 0;
        weight_mem[16'h135E] <= 0;
        weight_mem[16'h135F] <= 0;
        weight_mem[16'h1360] <= 0;
        weight_mem[16'h1361] <= 0;
        weight_mem[16'h1362] <= 0;
        weight_mem[16'h1363] <= 0;
        weight_mem[16'h1364] <= 0;
        weight_mem[16'h1365] <= 0;
        weight_mem[16'h1366] <= 0;
        weight_mem[16'h1367] <= 0;
        weight_mem[16'h1368] <= 0;
        weight_mem[16'h1369] <= 0;
        weight_mem[16'h136A] <= 0;
        weight_mem[16'h136B] <= 0;
        weight_mem[16'h136C] <= 0;
        weight_mem[16'h136D] <= 0;
        weight_mem[16'h136E] <= 0;
        weight_mem[16'h136F] <= 0;
        weight_mem[16'h1370] <= 0;
        weight_mem[16'h1371] <= 0;
        weight_mem[16'h1372] <= 0;
        weight_mem[16'h1373] <= 0;
        weight_mem[16'h1374] <= 0;
        weight_mem[16'h1375] <= 0;
        weight_mem[16'h1376] <= 0;
        weight_mem[16'h1377] <= 0;
        weight_mem[16'h1378] <= 0;
        weight_mem[16'h1379] <= 0;
        weight_mem[16'h137A] <= 0;
        weight_mem[16'h137B] <= 0;
        weight_mem[16'h137C] <= 0;
        weight_mem[16'h137D] <= 0;
        weight_mem[16'h137E] <= 0;
        weight_mem[16'h137F] <= 0;
        weight_mem[16'h1380] <= 0;
        weight_mem[16'h1381] <= 0;
        weight_mem[16'h1382] <= 0;
        weight_mem[16'h1383] <= 0;
        weight_mem[16'h1384] <= 0;
        weight_mem[16'h1385] <= 0;
        weight_mem[16'h1386] <= 0;
        weight_mem[16'h1387] <= 0;
        weight_mem[16'h1388] <= 0;
        weight_mem[16'h1389] <= 0;
        weight_mem[16'h138A] <= 0;
        weight_mem[16'h138B] <= 0;
        weight_mem[16'h138C] <= 0;
        weight_mem[16'h138D] <= 0;
        weight_mem[16'h138E] <= 0;
        weight_mem[16'h138F] <= 0;
        weight_mem[16'h1390] <= 0;
        weight_mem[16'h1391] <= 0;
        weight_mem[16'h1392] <= 0;
        weight_mem[16'h1393] <= 0;
        weight_mem[16'h1394] <= 0;
        weight_mem[16'h1395] <= 0;
        weight_mem[16'h1396] <= 0;
        weight_mem[16'h1397] <= 0;
        weight_mem[16'h1398] <= 0;
        weight_mem[16'h1399] <= 0;
        weight_mem[16'h139A] <= 0;
        weight_mem[16'h139B] <= 0;
        weight_mem[16'h139C] <= 0;
        weight_mem[16'h139D] <= 0;
        weight_mem[16'h139E] <= 0;
        weight_mem[16'h139F] <= 0;
        weight_mem[16'h13A0] <= 0;
        weight_mem[16'h13A1] <= 0;
        weight_mem[16'h13A2] <= 0;
        weight_mem[16'h13A3] <= 0;
        weight_mem[16'h13A4] <= 0;
        weight_mem[16'h13A5] <= 0;
        weight_mem[16'h13A6] <= 0;
        weight_mem[16'h13A7] <= 0;
        weight_mem[16'h13A8] <= 0;
        weight_mem[16'h13A9] <= 0;
        weight_mem[16'h13AA] <= 0;
        weight_mem[16'h13AB] <= 0;
        weight_mem[16'h13AC] <= 0;
        weight_mem[16'h13AD] <= 0;
        weight_mem[16'h13AE] <= 0;
        weight_mem[16'h13AF] <= 0;

        // layer 1 neuron 10
        weight_mem[16'h1400] <= 0;
        weight_mem[16'h1401] <= 0;
        weight_mem[16'h1402] <= 0;
        weight_mem[16'h1403] <= 0;
        weight_mem[16'h1404] <= 0;
        weight_mem[16'h1405] <= 0;
        weight_mem[16'h1406] <= 0;
        weight_mem[16'h1407] <= 0;
        weight_mem[16'h1408] <= 0;
        weight_mem[16'h1409] <= 0;
        weight_mem[16'h140A] <= 0;
        weight_mem[16'h140B] <= 0;
        weight_mem[16'h140C] <= 0;
        weight_mem[16'h140D] <= 0;
        weight_mem[16'h140E] <= 0;
        weight_mem[16'h140F] <= 0;
        weight_mem[16'h1410] <= 0;
        weight_mem[16'h1411] <= 0;
        weight_mem[16'h1412] <= 0;
        weight_mem[16'h1413] <= 0;
        weight_mem[16'h1414] <= 0;
        weight_mem[16'h1415] <= 0;
        weight_mem[16'h1416] <= 0;
        weight_mem[16'h1417] <= 0;
        weight_mem[16'h1418] <= 0;
        weight_mem[16'h1419] <= 0;
        weight_mem[16'h141A] <= 0;
        weight_mem[16'h141B] <= 0;
        weight_mem[16'h141C] <= 0;
        weight_mem[16'h141D] <= 0;
        weight_mem[16'h141E] <= 0;
        weight_mem[16'h141F] <= 0;
        weight_mem[16'h1420] <= 0;
        weight_mem[16'h1421] <= 0;
        weight_mem[16'h1422] <= 0;
        weight_mem[16'h1423] <= 0;
        weight_mem[16'h1424] <= 0;
        weight_mem[16'h1425] <= 0;
        weight_mem[16'h1426] <= 0;
        weight_mem[16'h1427] <= 0;
        weight_mem[16'h1428] <= 0;
        weight_mem[16'h1429] <= 0;
        weight_mem[16'h142A] <= 0;
        weight_mem[16'h142B] <= 0;
        weight_mem[16'h142C] <= 0;
        weight_mem[16'h142D] <= 0;
        weight_mem[16'h142E] <= 0;
        weight_mem[16'h142F] <= 0;
        weight_mem[16'h1430] <= 0;
        weight_mem[16'h1431] <= 0;
        weight_mem[16'h1432] <= 0;
        weight_mem[16'h1433] <= 0;
        weight_mem[16'h1434] <= 0;
        weight_mem[16'h1435] <= 0;
        weight_mem[16'h1436] <= 0;
        weight_mem[16'h1437] <= 0;
        weight_mem[16'h1438] <= 0;
        weight_mem[16'h1439] <= 0;
        weight_mem[16'h143A] <= 0;
        weight_mem[16'h143B] <= 0;
        weight_mem[16'h143C] <= 0;
        weight_mem[16'h143D] <= 0;
        weight_mem[16'h143E] <= 0;
        weight_mem[16'h143F] <= 0;
        weight_mem[16'h1440] <= 0;
        weight_mem[16'h1441] <= 0;
        weight_mem[16'h1442] <= 0;
        weight_mem[16'h1443] <= 0;
        weight_mem[16'h1444] <= 0;
        weight_mem[16'h1445] <= 0;
        weight_mem[16'h1446] <= 0;
        weight_mem[16'h1447] <= 0;
        weight_mem[16'h1448] <= 0;
        weight_mem[16'h1449] <= 0;
        weight_mem[16'h144A] <= 0;
        weight_mem[16'h144B] <= 0;
        weight_mem[16'h144C] <= 0;
        weight_mem[16'h144D] <= 0;
        weight_mem[16'h144E] <= 0;
        weight_mem[16'h144F] <= 0;
        weight_mem[16'h1450] <= 0;
        weight_mem[16'h1451] <= 0;
        weight_mem[16'h1452] <= 0;
        weight_mem[16'h1453] <= 0;
        weight_mem[16'h1454] <= 0;
        weight_mem[16'h1455] <= 0;
        weight_mem[16'h1456] <= 0;
        weight_mem[16'h1457] <= 0;
        weight_mem[16'h1458] <= 0;
        weight_mem[16'h1459] <= 0;
        weight_mem[16'h145A] <= 0;
        weight_mem[16'h145B] <= 0;
        weight_mem[16'h145C] <= 0;
        weight_mem[16'h145D] <= 0;
        weight_mem[16'h145E] <= 0;
        weight_mem[16'h145F] <= 0;
        weight_mem[16'h1460] <= 0;
        weight_mem[16'h1461] <= 0;
        weight_mem[16'h1462] <= 0;
        weight_mem[16'h1463] <= 0;
        weight_mem[16'h1464] <= 0;
        weight_mem[16'h1465] <= 0;
        weight_mem[16'h1466] <= 0;
        weight_mem[16'h1467] <= 0;
        weight_mem[16'h1468] <= 0;
        weight_mem[16'h1469] <= 0;
        weight_mem[16'h146A] <= 0;
        weight_mem[16'h146B] <= 0;
        weight_mem[16'h146C] <= 0;
        weight_mem[16'h146D] <= 0;
        weight_mem[16'h146E] <= 0;
        weight_mem[16'h146F] <= 0;
        weight_mem[16'h1470] <= 0;
        weight_mem[16'h1471] <= 0;
        weight_mem[16'h1472] <= 0;
        weight_mem[16'h1473] <= 0;
        weight_mem[16'h1474] <= 0;
        weight_mem[16'h1475] <= 0;
        weight_mem[16'h1476] <= 0;
        weight_mem[16'h1477] <= 0;
        weight_mem[16'h1478] <= 0;
        weight_mem[16'h1479] <= 0;
        weight_mem[16'h147A] <= 0;
        weight_mem[16'h147B] <= 0;
        weight_mem[16'h147C] <= 0;
        weight_mem[16'h147D] <= 0;
        weight_mem[16'h147E] <= 0;
        weight_mem[16'h147F] <= 0;
        weight_mem[16'h1480] <= 0;
        weight_mem[16'h1481] <= 0;
        weight_mem[16'h1482] <= 0;
        weight_mem[16'h1483] <= 0;
        weight_mem[16'h1484] <= 0;
        weight_mem[16'h1485] <= 0;
        weight_mem[16'h1486] <= 0;
        weight_mem[16'h1487] <= 0;
        weight_mem[16'h1488] <= 0;
        weight_mem[16'h1489] <= 0;
        weight_mem[16'h148A] <= 0;
        weight_mem[16'h148B] <= 0;
        weight_mem[16'h148C] <= 0;
        weight_mem[16'h148D] <= 0;
        weight_mem[16'h148E] <= 0;
        weight_mem[16'h148F] <= 0;
        weight_mem[16'h1490] <= 0;
        weight_mem[16'h1491] <= 0;
        weight_mem[16'h1492] <= 0;
        weight_mem[16'h1493] <= 0;
        weight_mem[16'h1494] <= 0;
        weight_mem[16'h1495] <= 0;
        weight_mem[16'h1496] <= 0;
        weight_mem[16'h1497] <= 0;
        weight_mem[16'h1498] <= 0;
        weight_mem[16'h1499] <= 0;
        weight_mem[16'h149A] <= 0;
        weight_mem[16'h149B] <= 0;
        weight_mem[16'h149C] <= 0;
        weight_mem[16'h149D] <= 0;
        weight_mem[16'h149E] <= 0;
        weight_mem[16'h149F] <= 0;
        weight_mem[16'h14A0] <= 0;
        weight_mem[16'h14A1] <= 0;
        weight_mem[16'h14A2] <= 0;
        weight_mem[16'h14A3] <= 0;
        weight_mem[16'h14A4] <= 0;
        weight_mem[16'h14A5] <= 0;
        weight_mem[16'h14A6] <= 0;
        weight_mem[16'h14A7] <= 0;
        weight_mem[16'h14A8] <= 0;
        weight_mem[16'h14A9] <= 0;
        weight_mem[16'h14AA] <= 0;
        weight_mem[16'h14AB] <= 0;
        weight_mem[16'h14AC] <= 0;
        weight_mem[16'h14AD] <= 0;
        weight_mem[16'h14AE] <= 0;
        weight_mem[16'h14AF] <= 0;
        weight_mem[16'h14B0] <= 0;
        weight_mem[16'h14B1] <= 0;
        weight_mem[16'h14B2] <= 0;
        weight_mem[16'h14B3] <= 0;
        weight_mem[16'h14B4] <= 0;
        weight_mem[16'h14B5] <= 0;
        weight_mem[16'h14B6] <= 0;
        weight_mem[16'h14B7] <= 0;
        weight_mem[16'h14B8] <= 0;
        weight_mem[16'h14B9] <= 0;
        weight_mem[16'h14BA] <= 0;
        weight_mem[16'h14BB] <= 0;
        weight_mem[16'h14BC] <= 0;
        weight_mem[16'h14BD] <= 0;
        weight_mem[16'h14BE] <= 0;
        weight_mem[16'h14BF] <= 0;
        weight_mem[16'h14C0] <= 0;
        weight_mem[16'h14C1] <= 0;
        weight_mem[16'h14C2] <= 0;
        weight_mem[16'h14C3] <= 0;
        weight_mem[16'h14C4] <= 0;
        weight_mem[16'h14C5] <= 0;
        weight_mem[16'h14C6] <= 0;
        weight_mem[16'h14C7] <= 0;
        weight_mem[16'h14C8] <= 0;
        weight_mem[16'h14C9] <= 0;
        weight_mem[16'h14CA] <= 0;
        weight_mem[16'h14CB] <= 0;
        weight_mem[16'h14CC] <= 0;
        weight_mem[16'h14CD] <= 0;
        weight_mem[16'h14CE] <= 0;
        weight_mem[16'h14CF] <= 0;
        weight_mem[16'h14D0] <= 0;
        weight_mem[16'h14D1] <= 0;
        weight_mem[16'h14D2] <= 0;
        weight_mem[16'h14D3] <= 0;
        weight_mem[16'h14D4] <= 0;
        weight_mem[16'h14D5] <= 0;
        weight_mem[16'h14D6] <= 0;
        weight_mem[16'h14D7] <= 0;
        weight_mem[16'h14D8] <= 0;
        weight_mem[16'h14D9] <= 0;
        weight_mem[16'h14DA] <= 0;
        weight_mem[16'h14DB] <= 0;
        weight_mem[16'h14DC] <= 0;
        weight_mem[16'h14DD] <= 0;
        weight_mem[16'h14DE] <= 0;
        weight_mem[16'h14DF] <= 0;
        weight_mem[16'h14E0] <= 0;
        weight_mem[16'h14E1] <= 0;
        weight_mem[16'h14E2] <= 0;
        weight_mem[16'h14E3] <= 0;
        weight_mem[16'h14E4] <= 0;
        weight_mem[16'h14E5] <= 0;
        weight_mem[16'h14E6] <= 0;
        weight_mem[16'h14E7] <= 0;
        weight_mem[16'h14E8] <= 0;
        weight_mem[16'h14E9] <= 0;
        weight_mem[16'h14EA] <= 0;
        weight_mem[16'h14EB] <= 0;
        weight_mem[16'h14EC] <= 0;
        weight_mem[16'h14ED] <= 0;
        weight_mem[16'h14EE] <= 0;
        weight_mem[16'h14EF] <= 0;
        weight_mem[16'h14F0] <= 0;
        weight_mem[16'h14F1] <= 0;
        weight_mem[16'h14F2] <= 0;
        weight_mem[16'h14F3] <= 0;
        weight_mem[16'h14F4] <= 0;
        weight_mem[16'h14F5] <= 0;
        weight_mem[16'h14F6] <= 0;
        weight_mem[16'h14F7] <= 0;
        weight_mem[16'h14F8] <= 0;
        weight_mem[16'h14F9] <= 0;
        weight_mem[16'h14FA] <= 0;
        weight_mem[16'h14FB] <= 0;
        weight_mem[16'h14FC] <= 0;
        weight_mem[16'h14FD] <= 0;
        weight_mem[16'h14FE] <= 0;
        weight_mem[16'h14FF] <= 0;
        weight_mem[16'h1500] <= 0;
        weight_mem[16'h1501] <= 0;
        weight_mem[16'h1502] <= 0;
        weight_mem[16'h1503] <= 0;
        weight_mem[16'h1504] <= 0;
        weight_mem[16'h1505] <= 0;
        weight_mem[16'h1506] <= 0;
        weight_mem[16'h1507] <= 0;
        weight_mem[16'h1508] <= 0;
        weight_mem[16'h1509] <= 0;
        weight_mem[16'h150A] <= 0;
        weight_mem[16'h150B] <= 0;
        weight_mem[16'h150C] <= 0;
        weight_mem[16'h150D] <= 0;
        weight_mem[16'h150E] <= 0;
        weight_mem[16'h150F] <= 0;
        weight_mem[16'h1510] <= 0;
        weight_mem[16'h1511] <= 0;
        weight_mem[16'h1512] <= 0;
        weight_mem[16'h1513] <= 0;
        weight_mem[16'h1514] <= 0;
        weight_mem[16'h1515] <= 0;
        weight_mem[16'h1516] <= 0;
        weight_mem[16'h1517] <= 0;
        weight_mem[16'h1518] <= 0;
        weight_mem[16'h1519] <= 0;
        weight_mem[16'h151A] <= 0;
        weight_mem[16'h151B] <= 0;
        weight_mem[16'h151C] <= 0;
        weight_mem[16'h151D] <= 0;
        weight_mem[16'h151E] <= 0;
        weight_mem[16'h151F] <= 0;
        weight_mem[16'h1520] <= 0;
        weight_mem[16'h1521] <= 0;
        weight_mem[16'h1522] <= 0;
        weight_mem[16'h1523] <= 0;
        weight_mem[16'h1524] <= 0;
        weight_mem[16'h1525] <= 0;
        weight_mem[16'h1526] <= 0;
        weight_mem[16'h1527] <= 0;
        weight_mem[16'h1528] <= 0;
        weight_mem[16'h1529] <= 0;
        weight_mem[16'h152A] <= 0;
        weight_mem[16'h152B] <= 0;
        weight_mem[16'h152C] <= 0;
        weight_mem[16'h152D] <= 0;
        weight_mem[16'h152E] <= 0;
        weight_mem[16'h152F] <= 0;
        weight_mem[16'h1530] <= 0;
        weight_mem[16'h1531] <= 0;
        weight_mem[16'h1532] <= 0;
        weight_mem[16'h1533] <= 0;
        weight_mem[16'h1534] <= 0;
        weight_mem[16'h1535] <= 0;
        weight_mem[16'h1536] <= 0;
        weight_mem[16'h1537] <= 0;
        weight_mem[16'h1538] <= 0;
        weight_mem[16'h1539] <= 0;
        weight_mem[16'h153A] <= 0;
        weight_mem[16'h153B] <= 0;
        weight_mem[16'h153C] <= 0;
        weight_mem[16'h153D] <= 0;
        weight_mem[16'h153E] <= 0;
        weight_mem[16'h153F] <= 0;
        weight_mem[16'h1540] <= 0;
        weight_mem[16'h1541] <= 0;
        weight_mem[16'h1542] <= 0;
        weight_mem[16'h1543] <= 0;
        weight_mem[16'h1544] <= 0;
        weight_mem[16'h1545] <= 0;
        weight_mem[16'h1546] <= 0;
        weight_mem[16'h1547] <= 0;
        weight_mem[16'h1548] <= 0;
        weight_mem[16'h1549] <= 0;
        weight_mem[16'h154A] <= 0;
        weight_mem[16'h154B] <= 0;
        weight_mem[16'h154C] <= 0;
        weight_mem[16'h154D] <= 0;
        weight_mem[16'h154E] <= 0;
        weight_mem[16'h154F] <= 0;
        weight_mem[16'h1550] <= 0;
        weight_mem[16'h1551] <= 0;
        weight_mem[16'h1552] <= 0;
        weight_mem[16'h1553] <= 0;
        weight_mem[16'h1554] <= 0;
        weight_mem[16'h1555] <= 0;
        weight_mem[16'h1556] <= 0;
        weight_mem[16'h1557] <= 0;
        weight_mem[16'h1558] <= 0;
        weight_mem[16'h1559] <= 0;
        weight_mem[16'h155A] <= 0;
        weight_mem[16'h155B] <= 0;
        weight_mem[16'h155C] <= 0;
        weight_mem[16'h155D] <= 0;
        weight_mem[16'h155E] <= 0;
        weight_mem[16'h155F] <= 0;
        weight_mem[16'h1560] <= 0;
        weight_mem[16'h1561] <= 0;
        weight_mem[16'h1562] <= 0;
        weight_mem[16'h1563] <= 0;
        weight_mem[16'h1564] <= 0;
        weight_mem[16'h1565] <= 0;
        weight_mem[16'h1566] <= 0;
        weight_mem[16'h1567] <= 0;
        weight_mem[16'h1568] <= 0;
        weight_mem[16'h1569] <= 0;
        weight_mem[16'h156A] <= 0;
        weight_mem[16'h156B] <= 0;
        weight_mem[16'h156C] <= 0;
        weight_mem[16'h156D] <= 0;
        weight_mem[16'h156E] <= 0;
        weight_mem[16'h156F] <= 0;
        weight_mem[16'h1570] <= 0;
        weight_mem[16'h1571] <= 0;
        weight_mem[16'h1572] <= 0;
        weight_mem[16'h1573] <= 0;
        weight_mem[16'h1574] <= 0;
        weight_mem[16'h1575] <= 0;
        weight_mem[16'h1576] <= 0;
        weight_mem[16'h1577] <= 0;
        weight_mem[16'h1578] <= 0;
        weight_mem[16'h1579] <= 0;
        weight_mem[16'h157A] <= 0;
        weight_mem[16'h157B] <= 0;
        weight_mem[16'h157C] <= 0;
        weight_mem[16'h157D] <= 0;
        weight_mem[16'h157E] <= 0;
        weight_mem[16'h157F] <= 0;
        weight_mem[16'h1580] <= 0;
        weight_mem[16'h1581] <= 0;
        weight_mem[16'h1582] <= 0;
        weight_mem[16'h1583] <= 0;
        weight_mem[16'h1584] <= 0;
        weight_mem[16'h1585] <= 0;
        weight_mem[16'h1586] <= 0;
        weight_mem[16'h1587] <= 0;
        weight_mem[16'h1588] <= 0;
        weight_mem[16'h1589] <= 0;
        weight_mem[16'h158A] <= 0;
        weight_mem[16'h158B] <= 0;
        weight_mem[16'h158C] <= 0;
        weight_mem[16'h158D] <= 0;
        weight_mem[16'h158E] <= 0;
        weight_mem[16'h158F] <= 0;
        weight_mem[16'h1590] <= 0;
        weight_mem[16'h1591] <= 0;
        weight_mem[16'h1592] <= 0;
        weight_mem[16'h1593] <= 0;
        weight_mem[16'h1594] <= 0;
        weight_mem[16'h1595] <= 0;
        weight_mem[16'h1596] <= 0;
        weight_mem[16'h1597] <= 0;
        weight_mem[16'h1598] <= 0;
        weight_mem[16'h1599] <= 0;
        weight_mem[16'h159A] <= 0;
        weight_mem[16'h159B] <= 0;
        weight_mem[16'h159C] <= 0;
        weight_mem[16'h159D] <= 0;
        weight_mem[16'h159E] <= 0;
        weight_mem[16'h159F] <= 0;
        weight_mem[16'h15A0] <= 0;
        weight_mem[16'h15A1] <= 0;
        weight_mem[16'h15A2] <= 0;
        weight_mem[16'h15A3] <= 0;
        weight_mem[16'h15A4] <= 0;
        weight_mem[16'h15A5] <= 0;
        weight_mem[16'h15A6] <= 0;
        weight_mem[16'h15A7] <= 0;
        weight_mem[16'h15A8] <= 0;
        weight_mem[16'h15A9] <= 0;
        weight_mem[16'h15AA] <= 0;
        weight_mem[16'h15AB] <= 0;
        weight_mem[16'h15AC] <= 0;
        weight_mem[16'h15AD] <= 0;
        weight_mem[16'h15AE] <= 0;
        weight_mem[16'h15AF] <= 0;

        // layer 1 neuron 11
        weight_mem[16'h1600] <= 0;
        weight_mem[16'h1601] <= 0;
        weight_mem[16'h1602] <= 0;
        weight_mem[16'h1603] <= 0;
        weight_mem[16'h1604] <= 0;
        weight_mem[16'h1605] <= 0;
        weight_mem[16'h1606] <= 0;
        weight_mem[16'h1607] <= 0;
        weight_mem[16'h1608] <= 0;
        weight_mem[16'h1609] <= 0;
        weight_mem[16'h160A] <= 0;
        weight_mem[16'h160B] <= 0;
        weight_mem[16'h160C] <= 0;
        weight_mem[16'h160D] <= 0;
        weight_mem[16'h160E] <= 0;
        weight_mem[16'h160F] <= 0;
        weight_mem[16'h1610] <= 0;
        weight_mem[16'h1611] <= 0;
        weight_mem[16'h1612] <= 0;
        weight_mem[16'h1613] <= 0;
        weight_mem[16'h1614] <= 0;
        weight_mem[16'h1615] <= 0;
        weight_mem[16'h1616] <= 0;
        weight_mem[16'h1617] <= 0;
        weight_mem[16'h1618] <= 0;
        weight_mem[16'h1619] <= 0;
        weight_mem[16'h161A] <= 0;
        weight_mem[16'h161B] <= 0;
        weight_mem[16'h161C] <= 0;
        weight_mem[16'h161D] <= 0;
        weight_mem[16'h161E] <= 0;
        weight_mem[16'h161F] <= 0;
        weight_mem[16'h1620] <= 0;
        weight_mem[16'h1621] <= 0;
        weight_mem[16'h1622] <= 0;
        weight_mem[16'h1623] <= 0;
        weight_mem[16'h1624] <= 0;
        weight_mem[16'h1625] <= 0;
        weight_mem[16'h1626] <= 0;
        weight_mem[16'h1627] <= 0;
        weight_mem[16'h1628] <= 0;
        weight_mem[16'h1629] <= 0;
        weight_mem[16'h162A] <= 0;
        weight_mem[16'h162B] <= 0;
        weight_mem[16'h162C] <= 0;
        weight_mem[16'h162D] <= 0;
        weight_mem[16'h162E] <= 0;
        weight_mem[16'h162F] <= 0;
        weight_mem[16'h1630] <= 0;
        weight_mem[16'h1631] <= 0;
        weight_mem[16'h1632] <= 0;
        weight_mem[16'h1633] <= 0;
        weight_mem[16'h1634] <= 0;
        weight_mem[16'h1635] <= 0;
        weight_mem[16'h1636] <= 0;
        weight_mem[16'h1637] <= 0;
        weight_mem[16'h1638] <= 0;
        weight_mem[16'h1639] <= 0;
        weight_mem[16'h163A] <= 0;
        weight_mem[16'h163B] <= 0;
        weight_mem[16'h163C] <= 0;
        weight_mem[16'h163D] <= 0;
        weight_mem[16'h163E] <= 0;
        weight_mem[16'h163F] <= 0;
        weight_mem[16'h1640] <= 0;
        weight_mem[16'h1641] <= 0;
        weight_mem[16'h1642] <= 0;
        weight_mem[16'h1643] <= 0;
        weight_mem[16'h1644] <= 0;
        weight_mem[16'h1645] <= 0;
        weight_mem[16'h1646] <= 0;
        weight_mem[16'h1647] <= 0;
        weight_mem[16'h1648] <= 0;
        weight_mem[16'h1649] <= 0;
        weight_mem[16'h164A] <= 0;
        weight_mem[16'h164B] <= 0;
        weight_mem[16'h164C] <= 0;
        weight_mem[16'h164D] <= 0;
        weight_mem[16'h164E] <= 0;
        weight_mem[16'h164F] <= 0;
        weight_mem[16'h1650] <= 0;
        weight_mem[16'h1651] <= 0;
        weight_mem[16'h1652] <= 0;
        weight_mem[16'h1653] <= 0;
        weight_mem[16'h1654] <= 0;
        weight_mem[16'h1655] <= 0;
        weight_mem[16'h1656] <= 0;
        weight_mem[16'h1657] <= 0;
        weight_mem[16'h1658] <= 0;
        weight_mem[16'h1659] <= 0;
        weight_mem[16'h165A] <= 0;
        weight_mem[16'h165B] <= 0;
        weight_mem[16'h165C] <= 0;
        weight_mem[16'h165D] <= 0;
        weight_mem[16'h165E] <= 0;
        weight_mem[16'h165F] <= 0;
        weight_mem[16'h1660] <= 0;
        weight_mem[16'h1661] <= 0;
        weight_mem[16'h1662] <= 0;
        weight_mem[16'h1663] <= 0;
        weight_mem[16'h1664] <= 0;
        weight_mem[16'h1665] <= 0;
        weight_mem[16'h1666] <= 0;
        weight_mem[16'h1667] <= 0;
        weight_mem[16'h1668] <= 0;
        weight_mem[16'h1669] <= 0;
        weight_mem[16'h166A] <= 0;
        weight_mem[16'h166B] <= 0;
        weight_mem[16'h166C] <= 0;
        weight_mem[16'h166D] <= 0;
        weight_mem[16'h166E] <= 0;
        weight_mem[16'h166F] <= 0;
        weight_mem[16'h1670] <= 0;
        weight_mem[16'h1671] <= 0;
        weight_mem[16'h1672] <= 0;
        weight_mem[16'h1673] <= 0;
        weight_mem[16'h1674] <= 0;
        weight_mem[16'h1675] <= 0;
        weight_mem[16'h1676] <= 0;
        weight_mem[16'h1677] <= 0;
        weight_mem[16'h1678] <= 0;
        weight_mem[16'h1679] <= 0;
        weight_mem[16'h167A] <= 0;
        weight_mem[16'h167B] <= 0;
        weight_mem[16'h167C] <= 0;
        weight_mem[16'h167D] <= 0;
        weight_mem[16'h167E] <= 0;
        weight_mem[16'h167F] <= 0;
        weight_mem[16'h1680] <= 0;
        weight_mem[16'h1681] <= 0;
        weight_mem[16'h1682] <= 0;
        weight_mem[16'h1683] <= 0;
        weight_mem[16'h1684] <= 0;
        weight_mem[16'h1685] <= 0;
        weight_mem[16'h1686] <= 0;
        weight_mem[16'h1687] <= 0;
        weight_mem[16'h1688] <= 0;
        weight_mem[16'h1689] <= 0;
        weight_mem[16'h168A] <= 0;
        weight_mem[16'h168B] <= 0;
        weight_mem[16'h168C] <= 0;
        weight_mem[16'h168D] <= 0;
        weight_mem[16'h168E] <= 0;
        weight_mem[16'h168F] <= 0;
        weight_mem[16'h1690] <= 0;
        weight_mem[16'h1691] <= 0;
        weight_mem[16'h1692] <= 0;
        weight_mem[16'h1693] <= 0;
        weight_mem[16'h1694] <= 0;
        weight_mem[16'h1695] <= 0;
        weight_mem[16'h1696] <= 0;
        weight_mem[16'h1697] <= 0;
        weight_mem[16'h1698] <= 0;
        weight_mem[16'h1699] <= 0;
        weight_mem[16'h169A] <= 0;
        weight_mem[16'h169B] <= 0;
        weight_mem[16'h169C] <= 0;
        weight_mem[16'h169D] <= 0;
        weight_mem[16'h169E] <= 0;
        weight_mem[16'h169F] <= 0;
        weight_mem[16'h16A0] <= 0;
        weight_mem[16'h16A1] <= 0;
        weight_mem[16'h16A2] <= 0;
        weight_mem[16'h16A3] <= 0;
        weight_mem[16'h16A4] <= 0;
        weight_mem[16'h16A5] <= 0;
        weight_mem[16'h16A6] <= 0;
        weight_mem[16'h16A7] <= 0;
        weight_mem[16'h16A8] <= 0;
        weight_mem[16'h16A9] <= 0;
        weight_mem[16'h16AA] <= 0;
        weight_mem[16'h16AB] <= 0;
        weight_mem[16'h16AC] <= 0;
        weight_mem[16'h16AD] <= 0;
        weight_mem[16'h16AE] <= 0;
        weight_mem[16'h16AF] <= 0;
        weight_mem[16'h16B0] <= 0;
        weight_mem[16'h16B1] <= 0;
        weight_mem[16'h16B2] <= 0;
        weight_mem[16'h16B3] <= 0;
        weight_mem[16'h16B4] <= 0;
        weight_mem[16'h16B5] <= 0;
        weight_mem[16'h16B6] <= 0;
        weight_mem[16'h16B7] <= 0;
        weight_mem[16'h16B8] <= 0;
        weight_mem[16'h16B9] <= 0;
        weight_mem[16'h16BA] <= 0;
        weight_mem[16'h16BB] <= 0;
        weight_mem[16'h16BC] <= 0;
        weight_mem[16'h16BD] <= 0;
        weight_mem[16'h16BE] <= 0;
        weight_mem[16'h16BF] <= 0;
        weight_mem[16'h16C0] <= 0;
        weight_mem[16'h16C1] <= 0;
        weight_mem[16'h16C2] <= 0;
        weight_mem[16'h16C3] <= 0;
        weight_mem[16'h16C4] <= 0;
        weight_mem[16'h16C5] <= 0;
        weight_mem[16'h16C6] <= 0;
        weight_mem[16'h16C7] <= 0;
        weight_mem[16'h16C8] <= 0;
        weight_mem[16'h16C9] <= 0;
        weight_mem[16'h16CA] <= 0;
        weight_mem[16'h16CB] <= 0;
        weight_mem[16'h16CC] <= 0;
        weight_mem[16'h16CD] <= 0;
        weight_mem[16'h16CE] <= 0;
        weight_mem[16'h16CF] <= 0;
        weight_mem[16'h16D0] <= 0;
        weight_mem[16'h16D1] <= 0;
        weight_mem[16'h16D2] <= 0;
        weight_mem[16'h16D3] <= 0;
        weight_mem[16'h16D4] <= 0;
        weight_mem[16'h16D5] <= 0;
        weight_mem[16'h16D6] <= 0;
        weight_mem[16'h16D7] <= 0;
        weight_mem[16'h16D8] <= 0;
        weight_mem[16'h16D9] <= 0;
        weight_mem[16'h16DA] <= 0;
        weight_mem[16'h16DB] <= 0;
        weight_mem[16'h16DC] <= 0;
        weight_mem[16'h16DD] <= 0;
        weight_mem[16'h16DE] <= 0;
        weight_mem[16'h16DF] <= 0;
        weight_mem[16'h16E0] <= 0;
        weight_mem[16'h16E1] <= 0;
        weight_mem[16'h16E2] <= 0;
        weight_mem[16'h16E3] <= 0;
        weight_mem[16'h16E4] <= 0;
        weight_mem[16'h16E5] <= 0;
        weight_mem[16'h16E6] <= 0;
        weight_mem[16'h16E7] <= 0;
        weight_mem[16'h16E8] <= 0;
        weight_mem[16'h16E9] <= 0;
        weight_mem[16'h16EA] <= 0;
        weight_mem[16'h16EB] <= 0;
        weight_mem[16'h16EC] <= 0;
        weight_mem[16'h16ED] <= 0;
        weight_mem[16'h16EE] <= 0;
        weight_mem[16'h16EF] <= 0;
        weight_mem[16'h16F0] <= 0;
        weight_mem[16'h16F1] <= 0;
        weight_mem[16'h16F2] <= 0;
        weight_mem[16'h16F3] <= 0;
        weight_mem[16'h16F4] <= 0;
        weight_mem[16'h16F5] <= 0;
        weight_mem[16'h16F6] <= 0;
        weight_mem[16'h16F7] <= 0;
        weight_mem[16'h16F8] <= 0;
        weight_mem[16'h16F9] <= 0;
        weight_mem[16'h16FA] <= 0;
        weight_mem[16'h16FB] <= 0;
        weight_mem[16'h16FC] <= 0;
        weight_mem[16'h16FD] <= 0;
        weight_mem[16'h16FE] <= 0;
        weight_mem[16'h16FF] <= 0;
        weight_mem[16'h1700] <= 0;
        weight_mem[16'h1701] <= 0;
        weight_mem[16'h1702] <= 0;
        weight_mem[16'h1703] <= 0;
        weight_mem[16'h1704] <= 0;
        weight_mem[16'h1705] <= 0;
        weight_mem[16'h1706] <= 0;
        weight_mem[16'h1707] <= 0;
        weight_mem[16'h1708] <= 0;
        weight_mem[16'h1709] <= 0;
        weight_mem[16'h170A] <= 0;
        weight_mem[16'h170B] <= 0;
        weight_mem[16'h170C] <= 0;
        weight_mem[16'h170D] <= 0;
        weight_mem[16'h170E] <= 0;
        weight_mem[16'h170F] <= 0;
        weight_mem[16'h1710] <= 0;
        weight_mem[16'h1711] <= 0;
        weight_mem[16'h1712] <= 0;
        weight_mem[16'h1713] <= 0;
        weight_mem[16'h1714] <= 0;
        weight_mem[16'h1715] <= 0;
        weight_mem[16'h1716] <= 0;
        weight_mem[16'h1717] <= 0;
        weight_mem[16'h1718] <= 0;
        weight_mem[16'h1719] <= 0;
        weight_mem[16'h171A] <= 0;
        weight_mem[16'h171B] <= 0;
        weight_mem[16'h171C] <= 0;
        weight_mem[16'h171D] <= 0;
        weight_mem[16'h171E] <= 0;
        weight_mem[16'h171F] <= 0;
        weight_mem[16'h1720] <= 0;
        weight_mem[16'h1721] <= 0;
        weight_mem[16'h1722] <= 0;
        weight_mem[16'h1723] <= 0;
        weight_mem[16'h1724] <= 0;
        weight_mem[16'h1725] <= 0;
        weight_mem[16'h1726] <= 0;
        weight_mem[16'h1727] <= 0;
        weight_mem[16'h1728] <= 0;
        weight_mem[16'h1729] <= 0;
        weight_mem[16'h172A] <= 0;
        weight_mem[16'h172B] <= 0;
        weight_mem[16'h172C] <= 0;
        weight_mem[16'h172D] <= 0;
        weight_mem[16'h172E] <= 0;
        weight_mem[16'h172F] <= 0;
        weight_mem[16'h1730] <= 0;
        weight_mem[16'h1731] <= 0;
        weight_mem[16'h1732] <= 0;
        weight_mem[16'h1733] <= 0;
        weight_mem[16'h1734] <= 0;
        weight_mem[16'h1735] <= 0;
        weight_mem[16'h1736] <= 0;
        weight_mem[16'h1737] <= 0;
        weight_mem[16'h1738] <= 0;
        weight_mem[16'h1739] <= 0;
        weight_mem[16'h173A] <= 0;
        weight_mem[16'h173B] <= 0;
        weight_mem[16'h173C] <= 0;
        weight_mem[16'h173D] <= 0;
        weight_mem[16'h173E] <= 0;
        weight_mem[16'h173F] <= 0;
        weight_mem[16'h1740] <= 0;
        weight_mem[16'h1741] <= 0;
        weight_mem[16'h1742] <= 0;
        weight_mem[16'h1743] <= 0;
        weight_mem[16'h1744] <= 0;
        weight_mem[16'h1745] <= 0;
        weight_mem[16'h1746] <= 0;
        weight_mem[16'h1747] <= 0;
        weight_mem[16'h1748] <= 0;
        weight_mem[16'h1749] <= 0;
        weight_mem[16'h174A] <= 0;
        weight_mem[16'h174B] <= 0;
        weight_mem[16'h174C] <= 0;
        weight_mem[16'h174D] <= 0;
        weight_mem[16'h174E] <= 0;
        weight_mem[16'h174F] <= 0;
        weight_mem[16'h1750] <= 0;
        weight_mem[16'h1751] <= 0;
        weight_mem[16'h1752] <= 0;
        weight_mem[16'h1753] <= 0;
        weight_mem[16'h1754] <= 0;
        weight_mem[16'h1755] <= 0;
        weight_mem[16'h1756] <= 0;
        weight_mem[16'h1757] <= 0;
        weight_mem[16'h1758] <= 0;
        weight_mem[16'h1759] <= 0;
        weight_mem[16'h175A] <= 0;
        weight_mem[16'h175B] <= 0;
        weight_mem[16'h175C] <= 0;
        weight_mem[16'h175D] <= 0;
        weight_mem[16'h175E] <= 0;
        weight_mem[16'h175F] <= 0;
        weight_mem[16'h1760] <= 0;
        weight_mem[16'h1761] <= 0;
        weight_mem[16'h1762] <= 0;
        weight_mem[16'h1763] <= 0;
        weight_mem[16'h1764] <= 0;
        weight_mem[16'h1765] <= 0;
        weight_mem[16'h1766] <= 0;
        weight_mem[16'h1767] <= 0;
        weight_mem[16'h1768] <= 0;
        weight_mem[16'h1769] <= 0;
        weight_mem[16'h176A] <= 0;
        weight_mem[16'h176B] <= 0;
        weight_mem[16'h176C] <= 0;
        weight_mem[16'h176D] <= 0;
        weight_mem[16'h176E] <= 0;
        weight_mem[16'h176F] <= 0;
        weight_mem[16'h1770] <= 0;
        weight_mem[16'h1771] <= 0;
        weight_mem[16'h1772] <= 0;
        weight_mem[16'h1773] <= 0;
        weight_mem[16'h1774] <= 0;
        weight_mem[16'h1775] <= 0;
        weight_mem[16'h1776] <= 0;
        weight_mem[16'h1777] <= 0;
        weight_mem[16'h1778] <= 0;
        weight_mem[16'h1779] <= 0;
        weight_mem[16'h177A] <= 0;
        weight_mem[16'h177B] <= 0;
        weight_mem[16'h177C] <= 0;
        weight_mem[16'h177D] <= 0;
        weight_mem[16'h177E] <= 0;
        weight_mem[16'h177F] <= 0;
        weight_mem[16'h1780] <= 0;
        weight_mem[16'h1781] <= 0;
        weight_mem[16'h1782] <= 0;
        weight_mem[16'h1783] <= 0;
        weight_mem[16'h1784] <= 0;
        weight_mem[16'h1785] <= 0;
        weight_mem[16'h1786] <= 0;
        weight_mem[16'h1787] <= 0;
        weight_mem[16'h1788] <= 0;
        weight_mem[16'h1789] <= 0;
        weight_mem[16'h178A] <= 0;
        weight_mem[16'h178B] <= 0;
        weight_mem[16'h178C] <= 0;
        weight_mem[16'h178D] <= 0;
        weight_mem[16'h178E] <= 0;
        weight_mem[16'h178F] <= 0;
        weight_mem[16'h1790] <= 0;
        weight_mem[16'h1791] <= 0;
        weight_mem[16'h1792] <= 0;
        weight_mem[16'h1793] <= 0;
        weight_mem[16'h1794] <= 0;
        weight_mem[16'h1795] <= 0;
        weight_mem[16'h1796] <= 0;
        weight_mem[16'h1797] <= 0;
        weight_mem[16'h1798] <= 0;
        weight_mem[16'h1799] <= 0;
        weight_mem[16'h179A] <= 0;
        weight_mem[16'h179B] <= 0;
        weight_mem[16'h179C] <= 0;
        weight_mem[16'h179D] <= 0;
        weight_mem[16'h179E] <= 0;
        weight_mem[16'h179F] <= 0;
        weight_mem[16'h17A0] <= 0;
        weight_mem[16'h17A1] <= 0;
        weight_mem[16'h17A2] <= 0;
        weight_mem[16'h17A3] <= 0;
        weight_mem[16'h17A4] <= 0;
        weight_mem[16'h17A5] <= 0;
        weight_mem[16'h17A6] <= 0;
        weight_mem[16'h17A7] <= 0;
        weight_mem[16'h17A8] <= 0;
        weight_mem[16'h17A9] <= 0;
        weight_mem[16'h17AA] <= 0;
        weight_mem[16'h17AB] <= 0;
        weight_mem[16'h17AC] <= 0;
        weight_mem[16'h17AD] <= 0;
        weight_mem[16'h17AE] <= 0;
        weight_mem[16'h17AF] <= 0;

        // layer 1 neuron 12
        weight_mem[16'h1800] <= 0;
        weight_mem[16'h1801] <= 0;
        weight_mem[16'h1802] <= 0;
        weight_mem[16'h1803] <= 0;
        weight_mem[16'h1804] <= 0;
        weight_mem[16'h1805] <= 0;
        weight_mem[16'h1806] <= 0;
        weight_mem[16'h1807] <= 0;
        weight_mem[16'h1808] <= 0;
        weight_mem[16'h1809] <= 0;
        weight_mem[16'h180A] <= 0;
        weight_mem[16'h180B] <= 0;
        weight_mem[16'h180C] <= 0;
        weight_mem[16'h180D] <= 0;
        weight_mem[16'h180E] <= 0;
        weight_mem[16'h180F] <= 0;
        weight_mem[16'h1810] <= 0;
        weight_mem[16'h1811] <= 0;
        weight_mem[16'h1812] <= 0;
        weight_mem[16'h1813] <= 0;
        weight_mem[16'h1814] <= 0;
        weight_mem[16'h1815] <= 0;
        weight_mem[16'h1816] <= 0;
        weight_mem[16'h1817] <= 0;
        weight_mem[16'h1818] <= 0;
        weight_mem[16'h1819] <= 0;
        weight_mem[16'h181A] <= 0;
        weight_mem[16'h181B] <= 0;
        weight_mem[16'h181C] <= 0;
        weight_mem[16'h181D] <= 0;
        weight_mem[16'h181E] <= 0;
        weight_mem[16'h181F] <= 0;
        weight_mem[16'h1820] <= 0;
        weight_mem[16'h1821] <= 0;
        weight_mem[16'h1822] <= 0;
        weight_mem[16'h1823] <= 0;
        weight_mem[16'h1824] <= 0;
        weight_mem[16'h1825] <= 0;
        weight_mem[16'h1826] <= 0;
        weight_mem[16'h1827] <= 0;
        weight_mem[16'h1828] <= 0;
        weight_mem[16'h1829] <= 0;
        weight_mem[16'h182A] <= 0;
        weight_mem[16'h182B] <= 0;
        weight_mem[16'h182C] <= 0;
        weight_mem[16'h182D] <= 0;
        weight_mem[16'h182E] <= 0;
        weight_mem[16'h182F] <= 0;
        weight_mem[16'h1830] <= 0;
        weight_mem[16'h1831] <= 0;
        weight_mem[16'h1832] <= 0;
        weight_mem[16'h1833] <= 0;
        weight_mem[16'h1834] <= 0;
        weight_mem[16'h1835] <= 0;
        weight_mem[16'h1836] <= 0;
        weight_mem[16'h1837] <= 0;
        weight_mem[16'h1838] <= 0;
        weight_mem[16'h1839] <= 0;
        weight_mem[16'h183A] <= 0;
        weight_mem[16'h183B] <= 0;
        weight_mem[16'h183C] <= 0;
        weight_mem[16'h183D] <= 0;
        weight_mem[16'h183E] <= 0;
        weight_mem[16'h183F] <= 0;
        weight_mem[16'h1840] <= 0;
        weight_mem[16'h1841] <= 0;
        weight_mem[16'h1842] <= 0;
        weight_mem[16'h1843] <= 0;
        weight_mem[16'h1844] <= 0;
        weight_mem[16'h1845] <= 0;
        weight_mem[16'h1846] <= 0;
        weight_mem[16'h1847] <= 0;
        weight_mem[16'h1848] <= 0;
        weight_mem[16'h1849] <= 0;
        weight_mem[16'h184A] <= 0;
        weight_mem[16'h184B] <= 0;
        weight_mem[16'h184C] <= 0;
        weight_mem[16'h184D] <= 0;
        weight_mem[16'h184E] <= 0;
        weight_mem[16'h184F] <= 0;
        weight_mem[16'h1850] <= 0;
        weight_mem[16'h1851] <= 0;
        weight_mem[16'h1852] <= 0;
        weight_mem[16'h1853] <= 0;
        weight_mem[16'h1854] <= 0;
        weight_mem[16'h1855] <= 0;
        weight_mem[16'h1856] <= 0;
        weight_mem[16'h1857] <= 0;
        weight_mem[16'h1858] <= 0;
        weight_mem[16'h1859] <= 0;
        weight_mem[16'h185A] <= 0;
        weight_mem[16'h185B] <= 0;
        weight_mem[16'h185C] <= 0;
        weight_mem[16'h185D] <= 0;
        weight_mem[16'h185E] <= 0;
        weight_mem[16'h185F] <= 0;
        weight_mem[16'h1860] <= 0;
        weight_mem[16'h1861] <= 0;
        weight_mem[16'h1862] <= 0;
        weight_mem[16'h1863] <= 0;
        weight_mem[16'h1864] <= 0;
        weight_mem[16'h1865] <= 0;
        weight_mem[16'h1866] <= 0;
        weight_mem[16'h1867] <= 0;
        weight_mem[16'h1868] <= 0;
        weight_mem[16'h1869] <= 0;
        weight_mem[16'h186A] <= 0;
        weight_mem[16'h186B] <= 0;
        weight_mem[16'h186C] <= 0;
        weight_mem[16'h186D] <= 0;
        weight_mem[16'h186E] <= 0;
        weight_mem[16'h186F] <= 0;
        weight_mem[16'h1870] <= 0;
        weight_mem[16'h1871] <= 0;
        weight_mem[16'h1872] <= 0;
        weight_mem[16'h1873] <= 0;
        weight_mem[16'h1874] <= 0;
        weight_mem[16'h1875] <= 0;
        weight_mem[16'h1876] <= 0;
        weight_mem[16'h1877] <= 0;
        weight_mem[16'h1878] <= 0;
        weight_mem[16'h1879] <= 0;
        weight_mem[16'h187A] <= 0;
        weight_mem[16'h187B] <= 0;
        weight_mem[16'h187C] <= 0;
        weight_mem[16'h187D] <= 0;
        weight_mem[16'h187E] <= 0;
        weight_mem[16'h187F] <= 0;
        weight_mem[16'h1880] <= 0;
        weight_mem[16'h1881] <= 0;
        weight_mem[16'h1882] <= 0;
        weight_mem[16'h1883] <= 0;
        weight_mem[16'h1884] <= 0;
        weight_mem[16'h1885] <= 0;
        weight_mem[16'h1886] <= 0;
        weight_mem[16'h1887] <= 0;
        weight_mem[16'h1888] <= 0;
        weight_mem[16'h1889] <= 0;
        weight_mem[16'h188A] <= 0;
        weight_mem[16'h188B] <= 0;
        weight_mem[16'h188C] <= 0;
        weight_mem[16'h188D] <= 0;
        weight_mem[16'h188E] <= 0;
        weight_mem[16'h188F] <= 0;
        weight_mem[16'h1890] <= 0;
        weight_mem[16'h1891] <= 0;
        weight_mem[16'h1892] <= 0;
        weight_mem[16'h1893] <= 0;
        weight_mem[16'h1894] <= 0;
        weight_mem[16'h1895] <= 0;
        weight_mem[16'h1896] <= 0;
        weight_mem[16'h1897] <= 0;
        weight_mem[16'h1898] <= 0;
        weight_mem[16'h1899] <= 0;
        weight_mem[16'h189A] <= 0;
        weight_mem[16'h189B] <= 0;
        weight_mem[16'h189C] <= 0;
        weight_mem[16'h189D] <= 0;
        weight_mem[16'h189E] <= 0;
        weight_mem[16'h189F] <= 0;
        weight_mem[16'h18A0] <= 0;
        weight_mem[16'h18A1] <= 0;
        weight_mem[16'h18A2] <= 0;
        weight_mem[16'h18A3] <= 0;
        weight_mem[16'h18A4] <= 0;
        weight_mem[16'h18A5] <= 0;
        weight_mem[16'h18A6] <= 0;
        weight_mem[16'h18A7] <= 0;
        weight_mem[16'h18A8] <= 0;
        weight_mem[16'h18A9] <= 0;
        weight_mem[16'h18AA] <= 0;
        weight_mem[16'h18AB] <= 0;
        weight_mem[16'h18AC] <= 0;
        weight_mem[16'h18AD] <= 0;
        weight_mem[16'h18AE] <= 0;
        weight_mem[16'h18AF] <= 0;
        weight_mem[16'h18B0] <= 0;
        weight_mem[16'h18B1] <= 0;
        weight_mem[16'h18B2] <= 0;
        weight_mem[16'h18B3] <= 0;
        weight_mem[16'h18B4] <= 0;
        weight_mem[16'h18B5] <= 0;
        weight_mem[16'h18B6] <= 0;
        weight_mem[16'h18B7] <= 0;
        weight_mem[16'h18B8] <= 0;
        weight_mem[16'h18B9] <= 0;
        weight_mem[16'h18BA] <= 0;
        weight_mem[16'h18BB] <= 0;
        weight_mem[16'h18BC] <= 0;
        weight_mem[16'h18BD] <= 0;
        weight_mem[16'h18BE] <= 0;
        weight_mem[16'h18BF] <= 0;
        weight_mem[16'h18C0] <= 0;
        weight_mem[16'h18C1] <= 0;
        weight_mem[16'h18C2] <= 0;
        weight_mem[16'h18C3] <= 0;
        weight_mem[16'h18C4] <= 0;
        weight_mem[16'h18C5] <= 0;
        weight_mem[16'h18C6] <= 0;
        weight_mem[16'h18C7] <= 0;
        weight_mem[16'h18C8] <= 0;
        weight_mem[16'h18C9] <= 0;
        weight_mem[16'h18CA] <= 0;
        weight_mem[16'h18CB] <= 0;
        weight_mem[16'h18CC] <= 0;
        weight_mem[16'h18CD] <= 0;
        weight_mem[16'h18CE] <= 0;
        weight_mem[16'h18CF] <= 0;
        weight_mem[16'h18D0] <= 0;
        weight_mem[16'h18D1] <= 0;
        weight_mem[16'h18D2] <= 0;
        weight_mem[16'h18D3] <= 0;
        weight_mem[16'h18D4] <= 0;
        weight_mem[16'h18D5] <= 0;
        weight_mem[16'h18D6] <= 0;
        weight_mem[16'h18D7] <= 0;
        weight_mem[16'h18D8] <= 0;
        weight_mem[16'h18D9] <= 0;
        weight_mem[16'h18DA] <= 0;
        weight_mem[16'h18DB] <= 0;
        weight_mem[16'h18DC] <= 0;
        weight_mem[16'h18DD] <= 0;
        weight_mem[16'h18DE] <= 0;
        weight_mem[16'h18DF] <= 0;
        weight_mem[16'h18E0] <= 0;
        weight_mem[16'h18E1] <= 0;
        weight_mem[16'h18E2] <= 0;
        weight_mem[16'h18E3] <= 0;
        weight_mem[16'h18E4] <= 0;
        weight_mem[16'h18E5] <= 0;
        weight_mem[16'h18E6] <= 0;
        weight_mem[16'h18E7] <= 0;
        weight_mem[16'h18E8] <= 0;
        weight_mem[16'h18E9] <= 0;
        weight_mem[16'h18EA] <= 0;
        weight_mem[16'h18EB] <= 0;
        weight_mem[16'h18EC] <= 0;
        weight_mem[16'h18ED] <= 0;
        weight_mem[16'h18EE] <= 0;
        weight_mem[16'h18EF] <= 0;
        weight_mem[16'h18F0] <= 0;
        weight_mem[16'h18F1] <= 0;
        weight_mem[16'h18F2] <= 0;
        weight_mem[16'h18F3] <= 0;
        weight_mem[16'h18F4] <= 0;
        weight_mem[16'h18F5] <= 0;
        weight_mem[16'h18F6] <= 0;
        weight_mem[16'h18F7] <= 0;
        weight_mem[16'h18F8] <= 0;
        weight_mem[16'h18F9] <= 0;
        weight_mem[16'h18FA] <= 0;
        weight_mem[16'h18FB] <= 0;
        weight_mem[16'h18FC] <= 0;
        weight_mem[16'h18FD] <= 0;
        weight_mem[16'h18FE] <= 0;
        weight_mem[16'h18FF] <= 0;
        weight_mem[16'h1900] <= 0;
        weight_mem[16'h1901] <= 0;
        weight_mem[16'h1902] <= 0;
        weight_mem[16'h1903] <= 0;
        weight_mem[16'h1904] <= 0;
        weight_mem[16'h1905] <= 0;
        weight_mem[16'h1906] <= 0;
        weight_mem[16'h1907] <= 0;
        weight_mem[16'h1908] <= 0;
        weight_mem[16'h1909] <= 0;
        weight_mem[16'h190A] <= 0;
        weight_mem[16'h190B] <= 0;
        weight_mem[16'h190C] <= 0;
        weight_mem[16'h190D] <= 0;
        weight_mem[16'h190E] <= 0;
        weight_mem[16'h190F] <= 0;
        weight_mem[16'h1910] <= 0;
        weight_mem[16'h1911] <= 0;
        weight_mem[16'h1912] <= 0;
        weight_mem[16'h1913] <= 0;
        weight_mem[16'h1914] <= 0;
        weight_mem[16'h1915] <= 0;
        weight_mem[16'h1916] <= 0;
        weight_mem[16'h1917] <= 0;
        weight_mem[16'h1918] <= 0;
        weight_mem[16'h1919] <= 0;
        weight_mem[16'h191A] <= 0;
        weight_mem[16'h191B] <= 0;
        weight_mem[16'h191C] <= 0;
        weight_mem[16'h191D] <= 0;
        weight_mem[16'h191E] <= 0;
        weight_mem[16'h191F] <= 0;
        weight_mem[16'h1920] <= 0;
        weight_mem[16'h1921] <= 0;
        weight_mem[16'h1922] <= 0;
        weight_mem[16'h1923] <= 0;
        weight_mem[16'h1924] <= 0;
        weight_mem[16'h1925] <= 0;
        weight_mem[16'h1926] <= 0;
        weight_mem[16'h1927] <= 0;
        weight_mem[16'h1928] <= 0;
        weight_mem[16'h1929] <= 0;
        weight_mem[16'h192A] <= 0;
        weight_mem[16'h192B] <= 0;
        weight_mem[16'h192C] <= 0;
        weight_mem[16'h192D] <= 0;
        weight_mem[16'h192E] <= 0;
        weight_mem[16'h192F] <= 0;
        weight_mem[16'h1930] <= 0;
        weight_mem[16'h1931] <= 0;
        weight_mem[16'h1932] <= 0;
        weight_mem[16'h1933] <= 0;
        weight_mem[16'h1934] <= 0;
        weight_mem[16'h1935] <= 0;
        weight_mem[16'h1936] <= 0;
        weight_mem[16'h1937] <= 0;
        weight_mem[16'h1938] <= 0;
        weight_mem[16'h1939] <= 0;
        weight_mem[16'h193A] <= 0;
        weight_mem[16'h193B] <= 0;
        weight_mem[16'h193C] <= 0;
        weight_mem[16'h193D] <= 0;
        weight_mem[16'h193E] <= 0;
        weight_mem[16'h193F] <= 0;
        weight_mem[16'h1940] <= 0;
        weight_mem[16'h1941] <= 0;
        weight_mem[16'h1942] <= 0;
        weight_mem[16'h1943] <= 0;
        weight_mem[16'h1944] <= 0;
        weight_mem[16'h1945] <= 0;
        weight_mem[16'h1946] <= 0;
        weight_mem[16'h1947] <= 0;
        weight_mem[16'h1948] <= 0;
        weight_mem[16'h1949] <= 0;
        weight_mem[16'h194A] <= 0;
        weight_mem[16'h194B] <= 0;
        weight_mem[16'h194C] <= 0;
        weight_mem[16'h194D] <= 0;
        weight_mem[16'h194E] <= 0;
        weight_mem[16'h194F] <= 0;
        weight_mem[16'h1950] <= 0;
        weight_mem[16'h1951] <= 0;
        weight_mem[16'h1952] <= 0;
        weight_mem[16'h1953] <= 0;
        weight_mem[16'h1954] <= 0;
        weight_mem[16'h1955] <= 0;
        weight_mem[16'h1956] <= 0;
        weight_mem[16'h1957] <= 0;
        weight_mem[16'h1958] <= 0;
        weight_mem[16'h1959] <= 0;
        weight_mem[16'h195A] <= 0;
        weight_mem[16'h195B] <= 0;
        weight_mem[16'h195C] <= 0;
        weight_mem[16'h195D] <= 0;
        weight_mem[16'h195E] <= 0;
        weight_mem[16'h195F] <= 0;
        weight_mem[16'h1960] <= 0;
        weight_mem[16'h1961] <= 0;
        weight_mem[16'h1962] <= 0;
        weight_mem[16'h1963] <= 0;
        weight_mem[16'h1964] <= 0;
        weight_mem[16'h1965] <= 0;
        weight_mem[16'h1966] <= 0;
        weight_mem[16'h1967] <= 0;
        weight_mem[16'h1968] <= 0;
        weight_mem[16'h1969] <= 0;
        weight_mem[16'h196A] <= 0;
        weight_mem[16'h196B] <= 0;
        weight_mem[16'h196C] <= 0;
        weight_mem[16'h196D] <= 0;
        weight_mem[16'h196E] <= 0;
        weight_mem[16'h196F] <= 0;
        weight_mem[16'h1970] <= 0;
        weight_mem[16'h1971] <= 0;
        weight_mem[16'h1972] <= 0;
        weight_mem[16'h1973] <= 0;
        weight_mem[16'h1974] <= 0;
        weight_mem[16'h1975] <= 0;
        weight_mem[16'h1976] <= 0;
        weight_mem[16'h1977] <= 0;
        weight_mem[16'h1978] <= 0;
        weight_mem[16'h1979] <= 0;
        weight_mem[16'h197A] <= 0;
        weight_mem[16'h197B] <= 0;
        weight_mem[16'h197C] <= 0;
        weight_mem[16'h197D] <= 0;
        weight_mem[16'h197E] <= 0;
        weight_mem[16'h197F] <= 0;
        weight_mem[16'h1980] <= 0;
        weight_mem[16'h1981] <= 0;
        weight_mem[16'h1982] <= 0;
        weight_mem[16'h1983] <= 0;
        weight_mem[16'h1984] <= 0;
        weight_mem[16'h1985] <= 0;
        weight_mem[16'h1986] <= 0;
        weight_mem[16'h1987] <= 0;
        weight_mem[16'h1988] <= 0;
        weight_mem[16'h1989] <= 0;
        weight_mem[16'h198A] <= 0;
        weight_mem[16'h198B] <= 0;
        weight_mem[16'h198C] <= 0;
        weight_mem[16'h198D] <= 0;
        weight_mem[16'h198E] <= 0;
        weight_mem[16'h198F] <= 0;
        weight_mem[16'h1990] <= 0;
        weight_mem[16'h1991] <= 0;
        weight_mem[16'h1992] <= 0;
        weight_mem[16'h1993] <= 0;
        weight_mem[16'h1994] <= 0;
        weight_mem[16'h1995] <= 0;
        weight_mem[16'h1996] <= 0;
        weight_mem[16'h1997] <= 0;
        weight_mem[16'h1998] <= 0;
        weight_mem[16'h1999] <= 0;
        weight_mem[16'h199A] <= 0;
        weight_mem[16'h199B] <= 0;
        weight_mem[16'h199C] <= 0;
        weight_mem[16'h199D] <= 0;
        weight_mem[16'h199E] <= 0;
        weight_mem[16'h199F] <= 0;
        weight_mem[16'h19A0] <= 0;
        weight_mem[16'h19A1] <= 0;
        weight_mem[16'h19A2] <= 0;
        weight_mem[16'h19A3] <= 0;
        weight_mem[16'h19A4] <= 0;
        weight_mem[16'h19A5] <= 0;
        weight_mem[16'h19A6] <= 0;
        weight_mem[16'h19A7] <= 0;
        weight_mem[16'h19A8] <= 0;
        weight_mem[16'h19A9] <= 0;
        weight_mem[16'h19AA] <= 0;
        weight_mem[16'h19AB] <= 0;
        weight_mem[16'h19AC] <= 0;
        weight_mem[16'h19AD] <= 0;
        weight_mem[16'h19AE] <= 0;
        weight_mem[16'h19AF] <= 0;

        // layer 1 neuron 13
        weight_mem[16'h1A00] <= 0;
        weight_mem[16'h1A01] <= 0;
        weight_mem[16'h1A02] <= 0;
        weight_mem[16'h1A03] <= 0;
        weight_mem[16'h1A04] <= 0;
        weight_mem[16'h1A05] <= 0;
        weight_mem[16'h1A06] <= 0;
        weight_mem[16'h1A07] <= 0;
        weight_mem[16'h1A08] <= 0;
        weight_mem[16'h1A09] <= 0;
        weight_mem[16'h1A0A] <= 0;
        weight_mem[16'h1A0B] <= 0;
        weight_mem[16'h1A0C] <= 0;
        weight_mem[16'h1A0D] <= 0;
        weight_mem[16'h1A0E] <= 0;
        weight_mem[16'h1A0F] <= 0;
        weight_mem[16'h1A10] <= 0;
        weight_mem[16'h1A11] <= 0;
        weight_mem[16'h1A12] <= 0;
        weight_mem[16'h1A13] <= 0;
        weight_mem[16'h1A14] <= 0;
        weight_mem[16'h1A15] <= 0;
        weight_mem[16'h1A16] <= 0;
        weight_mem[16'h1A17] <= 0;
        weight_mem[16'h1A18] <= 0;
        weight_mem[16'h1A19] <= 0;
        weight_mem[16'h1A1A] <= 0;
        weight_mem[16'h1A1B] <= 0;
        weight_mem[16'h1A1C] <= 0;
        weight_mem[16'h1A1D] <= 0;
        weight_mem[16'h1A1E] <= 0;
        weight_mem[16'h1A1F] <= 0;
        weight_mem[16'h1A20] <= 0;
        weight_mem[16'h1A21] <= 0;
        weight_mem[16'h1A22] <= 0;
        weight_mem[16'h1A23] <= 0;
        weight_mem[16'h1A24] <= 0;
        weight_mem[16'h1A25] <= 0;
        weight_mem[16'h1A26] <= 0;
        weight_mem[16'h1A27] <= 0;
        weight_mem[16'h1A28] <= 0;
        weight_mem[16'h1A29] <= 0;
        weight_mem[16'h1A2A] <= 0;
        weight_mem[16'h1A2B] <= 0;
        weight_mem[16'h1A2C] <= 0;
        weight_mem[16'h1A2D] <= 0;
        weight_mem[16'h1A2E] <= 0;
        weight_mem[16'h1A2F] <= 0;
        weight_mem[16'h1A30] <= 0;
        weight_mem[16'h1A31] <= 0;
        weight_mem[16'h1A32] <= 0;
        weight_mem[16'h1A33] <= 0;
        weight_mem[16'h1A34] <= 0;
        weight_mem[16'h1A35] <= 0;
        weight_mem[16'h1A36] <= 0;
        weight_mem[16'h1A37] <= 0;
        weight_mem[16'h1A38] <= 0;
        weight_mem[16'h1A39] <= 0;
        weight_mem[16'h1A3A] <= 0;
        weight_mem[16'h1A3B] <= 0;
        weight_mem[16'h1A3C] <= 0;
        weight_mem[16'h1A3D] <= 0;
        weight_mem[16'h1A3E] <= 0;
        weight_mem[16'h1A3F] <= 0;
        weight_mem[16'h1A40] <= 0;
        weight_mem[16'h1A41] <= 0;
        weight_mem[16'h1A42] <= 0;
        weight_mem[16'h1A43] <= 0;
        weight_mem[16'h1A44] <= 0;
        weight_mem[16'h1A45] <= 0;
        weight_mem[16'h1A46] <= 0;
        weight_mem[16'h1A47] <= 0;
        weight_mem[16'h1A48] <= 0;
        weight_mem[16'h1A49] <= 0;
        weight_mem[16'h1A4A] <= 0;
        weight_mem[16'h1A4B] <= 0;
        weight_mem[16'h1A4C] <= 0;
        weight_mem[16'h1A4D] <= 0;
        weight_mem[16'h1A4E] <= 0;
        weight_mem[16'h1A4F] <= 0;
        weight_mem[16'h1A50] <= 0;
        weight_mem[16'h1A51] <= 0;
        weight_mem[16'h1A52] <= 0;
        weight_mem[16'h1A53] <= 0;
        weight_mem[16'h1A54] <= 0;
        weight_mem[16'h1A55] <= 0;
        weight_mem[16'h1A56] <= 0;
        weight_mem[16'h1A57] <= 0;
        weight_mem[16'h1A58] <= 0;
        weight_mem[16'h1A59] <= 0;
        weight_mem[16'h1A5A] <= 0;
        weight_mem[16'h1A5B] <= 0;
        weight_mem[16'h1A5C] <= 0;
        weight_mem[16'h1A5D] <= 0;
        weight_mem[16'h1A5E] <= 0;
        weight_mem[16'h1A5F] <= 0;
        weight_mem[16'h1A60] <= 0;
        weight_mem[16'h1A61] <= 0;
        weight_mem[16'h1A62] <= 0;
        weight_mem[16'h1A63] <= 0;
        weight_mem[16'h1A64] <= 0;
        weight_mem[16'h1A65] <= 0;
        weight_mem[16'h1A66] <= 0;
        weight_mem[16'h1A67] <= 0;
        weight_mem[16'h1A68] <= 0;
        weight_mem[16'h1A69] <= 0;
        weight_mem[16'h1A6A] <= 0;
        weight_mem[16'h1A6B] <= 0;
        weight_mem[16'h1A6C] <= 0;
        weight_mem[16'h1A6D] <= 0;
        weight_mem[16'h1A6E] <= 0;
        weight_mem[16'h1A6F] <= 0;
        weight_mem[16'h1A70] <= 0;
        weight_mem[16'h1A71] <= 0;
        weight_mem[16'h1A72] <= 0;
        weight_mem[16'h1A73] <= 0;
        weight_mem[16'h1A74] <= 0;
        weight_mem[16'h1A75] <= 0;
        weight_mem[16'h1A76] <= 0;
        weight_mem[16'h1A77] <= 0;
        weight_mem[16'h1A78] <= 0;
        weight_mem[16'h1A79] <= 0;
        weight_mem[16'h1A7A] <= 0;
        weight_mem[16'h1A7B] <= 0;
        weight_mem[16'h1A7C] <= 0;
        weight_mem[16'h1A7D] <= 0;
        weight_mem[16'h1A7E] <= 0;
        weight_mem[16'h1A7F] <= 0;
        weight_mem[16'h1A80] <= 0;
        weight_mem[16'h1A81] <= 0;
        weight_mem[16'h1A82] <= 0;
        weight_mem[16'h1A83] <= 0;
        weight_mem[16'h1A84] <= 0;
        weight_mem[16'h1A85] <= 0;
        weight_mem[16'h1A86] <= 0;
        weight_mem[16'h1A87] <= 0;
        weight_mem[16'h1A88] <= 0;
        weight_mem[16'h1A89] <= 0;
        weight_mem[16'h1A8A] <= 0;
        weight_mem[16'h1A8B] <= 0;
        weight_mem[16'h1A8C] <= 0;
        weight_mem[16'h1A8D] <= 0;
        weight_mem[16'h1A8E] <= 0;
        weight_mem[16'h1A8F] <= 0;
        weight_mem[16'h1A90] <= 0;
        weight_mem[16'h1A91] <= 0;
        weight_mem[16'h1A92] <= 0;
        weight_mem[16'h1A93] <= 0;
        weight_mem[16'h1A94] <= 0;
        weight_mem[16'h1A95] <= 0;
        weight_mem[16'h1A96] <= 0;
        weight_mem[16'h1A97] <= 0;
        weight_mem[16'h1A98] <= 0;
        weight_mem[16'h1A99] <= 0;
        weight_mem[16'h1A9A] <= 0;
        weight_mem[16'h1A9B] <= 0;
        weight_mem[16'h1A9C] <= 0;
        weight_mem[16'h1A9D] <= 0;
        weight_mem[16'h1A9E] <= 0;
        weight_mem[16'h1A9F] <= 0;
        weight_mem[16'h1AA0] <= 0;
        weight_mem[16'h1AA1] <= 0;
        weight_mem[16'h1AA2] <= 0;
        weight_mem[16'h1AA3] <= 0;
        weight_mem[16'h1AA4] <= 0;
        weight_mem[16'h1AA5] <= 0;
        weight_mem[16'h1AA6] <= 0;
        weight_mem[16'h1AA7] <= 0;
        weight_mem[16'h1AA8] <= 0;
        weight_mem[16'h1AA9] <= 0;
        weight_mem[16'h1AAA] <= 0;
        weight_mem[16'h1AAB] <= 0;
        weight_mem[16'h1AAC] <= 0;
        weight_mem[16'h1AAD] <= 0;
        weight_mem[16'h1AAE] <= 0;
        weight_mem[16'h1AAF] <= 0;
        weight_mem[16'h1AB0] <= 0;
        weight_mem[16'h1AB1] <= 0;
        weight_mem[16'h1AB2] <= 0;
        weight_mem[16'h1AB3] <= 0;
        weight_mem[16'h1AB4] <= 0;
        weight_mem[16'h1AB5] <= 0;
        weight_mem[16'h1AB6] <= 0;
        weight_mem[16'h1AB7] <= 0;
        weight_mem[16'h1AB8] <= 0;
        weight_mem[16'h1AB9] <= 0;
        weight_mem[16'h1ABA] <= 0;
        weight_mem[16'h1ABB] <= 0;
        weight_mem[16'h1ABC] <= 0;
        weight_mem[16'h1ABD] <= 0;
        weight_mem[16'h1ABE] <= 0;
        weight_mem[16'h1ABF] <= 0;
        weight_mem[16'h1AC0] <= 0;
        weight_mem[16'h1AC1] <= 0;
        weight_mem[16'h1AC2] <= 0;
        weight_mem[16'h1AC3] <= 0;
        weight_mem[16'h1AC4] <= 0;
        weight_mem[16'h1AC5] <= 0;
        weight_mem[16'h1AC6] <= 0;
        weight_mem[16'h1AC7] <= 0;
        weight_mem[16'h1AC8] <= 0;
        weight_mem[16'h1AC9] <= 0;
        weight_mem[16'h1ACA] <= 0;
        weight_mem[16'h1ACB] <= 0;
        weight_mem[16'h1ACC] <= 0;
        weight_mem[16'h1ACD] <= 0;
        weight_mem[16'h1ACE] <= 0;
        weight_mem[16'h1ACF] <= 0;
        weight_mem[16'h1AD0] <= 0;
        weight_mem[16'h1AD1] <= 0;
        weight_mem[16'h1AD2] <= 0;
        weight_mem[16'h1AD3] <= 0;
        weight_mem[16'h1AD4] <= 0;
        weight_mem[16'h1AD5] <= 0;
        weight_mem[16'h1AD6] <= 0;
        weight_mem[16'h1AD7] <= 0;
        weight_mem[16'h1AD8] <= 0;
        weight_mem[16'h1AD9] <= 0;
        weight_mem[16'h1ADA] <= 0;
        weight_mem[16'h1ADB] <= 0;
        weight_mem[16'h1ADC] <= 0;
        weight_mem[16'h1ADD] <= 0;
        weight_mem[16'h1ADE] <= 0;
        weight_mem[16'h1ADF] <= 0;
        weight_mem[16'h1AE0] <= 0;
        weight_mem[16'h1AE1] <= 0;
        weight_mem[16'h1AE2] <= 0;
        weight_mem[16'h1AE3] <= 0;
        weight_mem[16'h1AE4] <= 0;
        weight_mem[16'h1AE5] <= 0;
        weight_mem[16'h1AE6] <= 0;
        weight_mem[16'h1AE7] <= 0;
        weight_mem[16'h1AE8] <= 0;
        weight_mem[16'h1AE9] <= 0;
        weight_mem[16'h1AEA] <= 0;
        weight_mem[16'h1AEB] <= 0;
        weight_mem[16'h1AEC] <= 0;
        weight_mem[16'h1AED] <= 0;
        weight_mem[16'h1AEE] <= 0;
        weight_mem[16'h1AEF] <= 0;
        weight_mem[16'h1AF0] <= 0;
        weight_mem[16'h1AF1] <= 0;
        weight_mem[16'h1AF2] <= 0;
        weight_mem[16'h1AF3] <= 0;
        weight_mem[16'h1AF4] <= 0;
        weight_mem[16'h1AF5] <= 0;
        weight_mem[16'h1AF6] <= 0;
        weight_mem[16'h1AF7] <= 0;
        weight_mem[16'h1AF8] <= 0;
        weight_mem[16'h1AF9] <= 0;
        weight_mem[16'h1AFA] <= 0;
        weight_mem[16'h1AFB] <= 0;
        weight_mem[16'h1AFC] <= 0;
        weight_mem[16'h1AFD] <= 0;
        weight_mem[16'h1AFE] <= 0;
        weight_mem[16'h1AFF] <= 0;
        weight_mem[16'h1B00] <= 0;
        weight_mem[16'h1B01] <= 0;
        weight_mem[16'h1B02] <= 0;
        weight_mem[16'h1B03] <= 0;
        weight_mem[16'h1B04] <= 0;
        weight_mem[16'h1B05] <= 0;
        weight_mem[16'h1B06] <= 0;
        weight_mem[16'h1B07] <= 0;
        weight_mem[16'h1B08] <= 0;
        weight_mem[16'h1B09] <= 0;
        weight_mem[16'h1B0A] <= 0;
        weight_mem[16'h1B0B] <= 0;
        weight_mem[16'h1B0C] <= 0;
        weight_mem[16'h1B0D] <= 0;
        weight_mem[16'h1B0E] <= 0;
        weight_mem[16'h1B0F] <= 0;
        weight_mem[16'h1B10] <= 0;
        weight_mem[16'h1B11] <= 0;
        weight_mem[16'h1B12] <= 0;
        weight_mem[16'h1B13] <= 0;
        weight_mem[16'h1B14] <= 0;
        weight_mem[16'h1B15] <= 0;
        weight_mem[16'h1B16] <= 0;
        weight_mem[16'h1B17] <= 0;
        weight_mem[16'h1B18] <= 0;
        weight_mem[16'h1B19] <= 0;
        weight_mem[16'h1B1A] <= 0;
        weight_mem[16'h1B1B] <= 0;
        weight_mem[16'h1B1C] <= 0;
        weight_mem[16'h1B1D] <= 0;
        weight_mem[16'h1B1E] <= 0;
        weight_mem[16'h1B1F] <= 0;
        weight_mem[16'h1B20] <= 0;
        weight_mem[16'h1B21] <= 0;
        weight_mem[16'h1B22] <= 0;
        weight_mem[16'h1B23] <= 0;
        weight_mem[16'h1B24] <= 0;
        weight_mem[16'h1B25] <= 0;
        weight_mem[16'h1B26] <= 0;
        weight_mem[16'h1B27] <= 0;
        weight_mem[16'h1B28] <= 0;
        weight_mem[16'h1B29] <= 0;
        weight_mem[16'h1B2A] <= 0;
        weight_mem[16'h1B2B] <= 0;
        weight_mem[16'h1B2C] <= 0;
        weight_mem[16'h1B2D] <= 0;
        weight_mem[16'h1B2E] <= 0;
        weight_mem[16'h1B2F] <= 0;
        weight_mem[16'h1B30] <= 0;
        weight_mem[16'h1B31] <= 0;
        weight_mem[16'h1B32] <= 0;
        weight_mem[16'h1B33] <= 0;
        weight_mem[16'h1B34] <= 0;
        weight_mem[16'h1B35] <= 0;
        weight_mem[16'h1B36] <= 0;
        weight_mem[16'h1B37] <= 0;
        weight_mem[16'h1B38] <= 0;
        weight_mem[16'h1B39] <= 0;
        weight_mem[16'h1B3A] <= 0;
        weight_mem[16'h1B3B] <= 0;
        weight_mem[16'h1B3C] <= 0;
        weight_mem[16'h1B3D] <= 0;
        weight_mem[16'h1B3E] <= 0;
        weight_mem[16'h1B3F] <= 0;
        weight_mem[16'h1B40] <= 0;
        weight_mem[16'h1B41] <= 0;
        weight_mem[16'h1B42] <= 0;
        weight_mem[16'h1B43] <= 0;
        weight_mem[16'h1B44] <= 0;
        weight_mem[16'h1B45] <= 0;
        weight_mem[16'h1B46] <= 0;
        weight_mem[16'h1B47] <= 0;
        weight_mem[16'h1B48] <= 0;
        weight_mem[16'h1B49] <= 0;
        weight_mem[16'h1B4A] <= 0;
        weight_mem[16'h1B4B] <= 0;
        weight_mem[16'h1B4C] <= 0;
        weight_mem[16'h1B4D] <= 0;
        weight_mem[16'h1B4E] <= 0;
        weight_mem[16'h1B4F] <= 0;
        weight_mem[16'h1B50] <= 0;
        weight_mem[16'h1B51] <= 0;
        weight_mem[16'h1B52] <= 0;
        weight_mem[16'h1B53] <= 0;
        weight_mem[16'h1B54] <= 0;
        weight_mem[16'h1B55] <= 0;
        weight_mem[16'h1B56] <= 0;
        weight_mem[16'h1B57] <= 0;
        weight_mem[16'h1B58] <= 0;
        weight_mem[16'h1B59] <= 0;
        weight_mem[16'h1B5A] <= 0;
        weight_mem[16'h1B5B] <= 0;
        weight_mem[16'h1B5C] <= 0;
        weight_mem[16'h1B5D] <= 0;
        weight_mem[16'h1B5E] <= 0;
        weight_mem[16'h1B5F] <= 0;
        weight_mem[16'h1B60] <= 0;
        weight_mem[16'h1B61] <= 0;
        weight_mem[16'h1B62] <= 0;
        weight_mem[16'h1B63] <= 0;
        weight_mem[16'h1B64] <= 0;
        weight_mem[16'h1B65] <= 0;
        weight_mem[16'h1B66] <= 0;
        weight_mem[16'h1B67] <= 0;
        weight_mem[16'h1B68] <= 0;
        weight_mem[16'h1B69] <= 0;
        weight_mem[16'h1B6A] <= 0;
        weight_mem[16'h1B6B] <= 0;
        weight_mem[16'h1B6C] <= 0;
        weight_mem[16'h1B6D] <= 0;
        weight_mem[16'h1B6E] <= 0;
        weight_mem[16'h1B6F] <= 0;
        weight_mem[16'h1B70] <= 0;
        weight_mem[16'h1B71] <= 0;
        weight_mem[16'h1B72] <= 0;
        weight_mem[16'h1B73] <= 0;
        weight_mem[16'h1B74] <= 0;
        weight_mem[16'h1B75] <= 0;
        weight_mem[16'h1B76] <= 0;
        weight_mem[16'h1B77] <= 0;
        weight_mem[16'h1B78] <= 0;
        weight_mem[16'h1B79] <= 0;
        weight_mem[16'h1B7A] <= 0;
        weight_mem[16'h1B7B] <= 0;
        weight_mem[16'h1B7C] <= 0;
        weight_mem[16'h1B7D] <= 0;
        weight_mem[16'h1B7E] <= 0;
        weight_mem[16'h1B7F] <= 0;
        weight_mem[16'h1B80] <= 0;
        weight_mem[16'h1B81] <= 0;
        weight_mem[16'h1B82] <= 0;
        weight_mem[16'h1B83] <= 0;
        weight_mem[16'h1B84] <= 0;
        weight_mem[16'h1B85] <= 0;
        weight_mem[16'h1B86] <= 0;
        weight_mem[16'h1B87] <= 0;
        weight_mem[16'h1B88] <= 0;
        weight_mem[16'h1B89] <= 0;
        weight_mem[16'h1B8A] <= 0;
        weight_mem[16'h1B8B] <= 0;
        weight_mem[16'h1B8C] <= 0;
        weight_mem[16'h1B8D] <= 0;
        weight_mem[16'h1B8E] <= 0;
        weight_mem[16'h1B8F] <= 0;
        weight_mem[16'h1B90] <= 0;
        weight_mem[16'h1B91] <= 0;
        weight_mem[16'h1B92] <= 0;
        weight_mem[16'h1B93] <= 0;
        weight_mem[16'h1B94] <= 0;
        weight_mem[16'h1B95] <= 0;
        weight_mem[16'h1B96] <= 0;
        weight_mem[16'h1B97] <= 0;
        weight_mem[16'h1B98] <= 0;
        weight_mem[16'h1B99] <= 0;
        weight_mem[16'h1B9A] <= 0;
        weight_mem[16'h1B9B] <= 0;
        weight_mem[16'h1B9C] <= 0;
        weight_mem[16'h1B9D] <= 0;
        weight_mem[16'h1B9E] <= 0;
        weight_mem[16'h1B9F] <= 0;
        weight_mem[16'h1BA0] <= 0;
        weight_mem[16'h1BA1] <= 0;
        weight_mem[16'h1BA2] <= 0;
        weight_mem[16'h1BA3] <= 0;
        weight_mem[16'h1BA4] <= 0;
        weight_mem[16'h1BA5] <= 0;
        weight_mem[16'h1BA6] <= 0;
        weight_mem[16'h1BA7] <= 0;
        weight_mem[16'h1BA8] <= 0;
        weight_mem[16'h1BA9] <= 0;
        weight_mem[16'h1BAA] <= 0;
        weight_mem[16'h1BAB] <= 0;
        weight_mem[16'h1BAC] <= 0;
        weight_mem[16'h1BAD] <= 0;
        weight_mem[16'h1BAE] <= 0;
        weight_mem[16'h1BAF] <= 0;

        // layer 1 neuron 14
        weight_mem[16'h1C00] <= 0;
        weight_mem[16'h1C01] <= 0;
        weight_mem[16'h1C02] <= 0;
        weight_mem[16'h1C03] <= 0;
        weight_mem[16'h1C04] <= 0;
        weight_mem[16'h1C05] <= 0;
        weight_mem[16'h1C06] <= 0;
        weight_mem[16'h1C07] <= 0;
        weight_mem[16'h1C08] <= 0;
        weight_mem[16'h1C09] <= 0;
        weight_mem[16'h1C0A] <= 0;
        weight_mem[16'h1C0B] <= 0;
        weight_mem[16'h1C0C] <= 0;
        weight_mem[16'h1C0D] <= 0;
        weight_mem[16'h1C0E] <= 0;
        weight_mem[16'h1C0F] <= 0;
        weight_mem[16'h1C10] <= 0;
        weight_mem[16'h1C11] <= 0;
        weight_mem[16'h1C12] <= 0;
        weight_mem[16'h1C13] <= 0;
        weight_mem[16'h1C14] <= 0;
        weight_mem[16'h1C15] <= 0;
        weight_mem[16'h1C16] <= 0;
        weight_mem[16'h1C17] <= 0;
        weight_mem[16'h1C18] <= 0;
        weight_mem[16'h1C19] <= 0;
        weight_mem[16'h1C1A] <= 0;
        weight_mem[16'h1C1B] <= 0;
        weight_mem[16'h1C1C] <= 0;
        weight_mem[16'h1C1D] <= 0;
        weight_mem[16'h1C1E] <= 0;
        weight_mem[16'h1C1F] <= 0;
        weight_mem[16'h1C20] <= 0;
        weight_mem[16'h1C21] <= 0;
        weight_mem[16'h1C22] <= 0;
        weight_mem[16'h1C23] <= 0;
        weight_mem[16'h1C24] <= 0;
        weight_mem[16'h1C25] <= 0;
        weight_mem[16'h1C26] <= 0;
        weight_mem[16'h1C27] <= 0;
        weight_mem[16'h1C28] <= 0;
        weight_mem[16'h1C29] <= 0;
        weight_mem[16'h1C2A] <= 0;
        weight_mem[16'h1C2B] <= 0;
        weight_mem[16'h1C2C] <= 0;
        weight_mem[16'h1C2D] <= 0;
        weight_mem[16'h1C2E] <= 0;
        weight_mem[16'h1C2F] <= 0;
        weight_mem[16'h1C30] <= 0;
        weight_mem[16'h1C31] <= 0;
        weight_mem[16'h1C32] <= 0;
        weight_mem[16'h1C33] <= 0;
        weight_mem[16'h1C34] <= 0;
        weight_mem[16'h1C35] <= 0;
        weight_mem[16'h1C36] <= 0;
        weight_mem[16'h1C37] <= 0;
        weight_mem[16'h1C38] <= 0;
        weight_mem[16'h1C39] <= 0;
        weight_mem[16'h1C3A] <= 0;
        weight_mem[16'h1C3B] <= 0;
        weight_mem[16'h1C3C] <= 0;
        weight_mem[16'h1C3D] <= 0;
        weight_mem[16'h1C3E] <= 0;
        weight_mem[16'h1C3F] <= 0;
        weight_mem[16'h1C40] <= 0;
        weight_mem[16'h1C41] <= 0;
        weight_mem[16'h1C42] <= 0;
        weight_mem[16'h1C43] <= 0;
        weight_mem[16'h1C44] <= 0;
        weight_mem[16'h1C45] <= 0;
        weight_mem[16'h1C46] <= 0;
        weight_mem[16'h1C47] <= 0;
        weight_mem[16'h1C48] <= 0;
        weight_mem[16'h1C49] <= 0;
        weight_mem[16'h1C4A] <= 0;
        weight_mem[16'h1C4B] <= 0;
        weight_mem[16'h1C4C] <= 0;
        weight_mem[16'h1C4D] <= 0;
        weight_mem[16'h1C4E] <= 0;
        weight_mem[16'h1C4F] <= 0;
        weight_mem[16'h1C50] <= 0;
        weight_mem[16'h1C51] <= 0;
        weight_mem[16'h1C52] <= 0;
        weight_mem[16'h1C53] <= 0;
        weight_mem[16'h1C54] <= 0;
        weight_mem[16'h1C55] <= 0;
        weight_mem[16'h1C56] <= 0;
        weight_mem[16'h1C57] <= 0;
        weight_mem[16'h1C58] <= 0;
        weight_mem[16'h1C59] <= 0;
        weight_mem[16'h1C5A] <= 0;
        weight_mem[16'h1C5B] <= 0;
        weight_mem[16'h1C5C] <= 0;
        weight_mem[16'h1C5D] <= 0;
        weight_mem[16'h1C5E] <= 0;
        weight_mem[16'h1C5F] <= 0;
        weight_mem[16'h1C60] <= 0;
        weight_mem[16'h1C61] <= 0;
        weight_mem[16'h1C62] <= 0;
        weight_mem[16'h1C63] <= 0;
        weight_mem[16'h1C64] <= 0;
        weight_mem[16'h1C65] <= 0;
        weight_mem[16'h1C66] <= 0;
        weight_mem[16'h1C67] <= 0;
        weight_mem[16'h1C68] <= 0;
        weight_mem[16'h1C69] <= 0;
        weight_mem[16'h1C6A] <= 0;
        weight_mem[16'h1C6B] <= 0;
        weight_mem[16'h1C6C] <= 0;
        weight_mem[16'h1C6D] <= 0;
        weight_mem[16'h1C6E] <= 0;
        weight_mem[16'h1C6F] <= 0;
        weight_mem[16'h1C70] <= 0;
        weight_mem[16'h1C71] <= 0;
        weight_mem[16'h1C72] <= 0;
        weight_mem[16'h1C73] <= 0;
        weight_mem[16'h1C74] <= 0;
        weight_mem[16'h1C75] <= 0;
        weight_mem[16'h1C76] <= 0;
        weight_mem[16'h1C77] <= 0;
        weight_mem[16'h1C78] <= 0;
        weight_mem[16'h1C79] <= 0;
        weight_mem[16'h1C7A] <= 0;
        weight_mem[16'h1C7B] <= 0;
        weight_mem[16'h1C7C] <= 0;
        weight_mem[16'h1C7D] <= 0;
        weight_mem[16'h1C7E] <= 0;
        weight_mem[16'h1C7F] <= 0;
        weight_mem[16'h1C80] <= 0;
        weight_mem[16'h1C81] <= 0;
        weight_mem[16'h1C82] <= 0;
        weight_mem[16'h1C83] <= 0;
        weight_mem[16'h1C84] <= 0;
        weight_mem[16'h1C85] <= 0;
        weight_mem[16'h1C86] <= 0;
        weight_mem[16'h1C87] <= 0;
        weight_mem[16'h1C88] <= 0;
        weight_mem[16'h1C89] <= 0;
        weight_mem[16'h1C8A] <= 0;
        weight_mem[16'h1C8B] <= 0;
        weight_mem[16'h1C8C] <= 0;
        weight_mem[16'h1C8D] <= 0;
        weight_mem[16'h1C8E] <= 0;
        weight_mem[16'h1C8F] <= 0;
        weight_mem[16'h1C90] <= 0;
        weight_mem[16'h1C91] <= 0;
        weight_mem[16'h1C92] <= 0;
        weight_mem[16'h1C93] <= 0;
        weight_mem[16'h1C94] <= 0;
        weight_mem[16'h1C95] <= 0;
        weight_mem[16'h1C96] <= 0;
        weight_mem[16'h1C97] <= 0;
        weight_mem[16'h1C98] <= 0;
        weight_mem[16'h1C99] <= 0;
        weight_mem[16'h1C9A] <= 0;
        weight_mem[16'h1C9B] <= 0;
        weight_mem[16'h1C9C] <= 0;
        weight_mem[16'h1C9D] <= 0;
        weight_mem[16'h1C9E] <= 0;
        weight_mem[16'h1C9F] <= 0;
        weight_mem[16'h1CA0] <= 0;
        weight_mem[16'h1CA1] <= 0;
        weight_mem[16'h1CA2] <= 0;
        weight_mem[16'h1CA3] <= 0;
        weight_mem[16'h1CA4] <= 0;
        weight_mem[16'h1CA5] <= 0;
        weight_mem[16'h1CA6] <= 0;
        weight_mem[16'h1CA7] <= 0;
        weight_mem[16'h1CA8] <= 0;
        weight_mem[16'h1CA9] <= 0;
        weight_mem[16'h1CAA] <= 0;
        weight_mem[16'h1CAB] <= 0;
        weight_mem[16'h1CAC] <= 0;
        weight_mem[16'h1CAD] <= 0;
        weight_mem[16'h1CAE] <= 0;
        weight_mem[16'h1CAF] <= 0;
        weight_mem[16'h1CB0] <= 0;
        weight_mem[16'h1CB1] <= 0;
        weight_mem[16'h1CB2] <= 0;
        weight_mem[16'h1CB3] <= 0;
        weight_mem[16'h1CB4] <= 0;
        weight_mem[16'h1CB5] <= 0;
        weight_mem[16'h1CB6] <= 0;
        weight_mem[16'h1CB7] <= 0;
        weight_mem[16'h1CB8] <= 0;
        weight_mem[16'h1CB9] <= 0;
        weight_mem[16'h1CBA] <= 0;
        weight_mem[16'h1CBB] <= 0;
        weight_mem[16'h1CBC] <= 0;
        weight_mem[16'h1CBD] <= 0;
        weight_mem[16'h1CBE] <= 0;
        weight_mem[16'h1CBF] <= 0;
        weight_mem[16'h1CC0] <= 0;
        weight_mem[16'h1CC1] <= 0;
        weight_mem[16'h1CC2] <= 0;
        weight_mem[16'h1CC3] <= 0;
        weight_mem[16'h1CC4] <= 0;
        weight_mem[16'h1CC5] <= 0;
        weight_mem[16'h1CC6] <= 0;
        weight_mem[16'h1CC7] <= 0;
        weight_mem[16'h1CC8] <= 0;
        weight_mem[16'h1CC9] <= 0;
        weight_mem[16'h1CCA] <= 0;
        weight_mem[16'h1CCB] <= 0;
        weight_mem[16'h1CCC] <= 0;
        weight_mem[16'h1CCD] <= 0;
        weight_mem[16'h1CCE] <= 0;
        weight_mem[16'h1CCF] <= 0;
        weight_mem[16'h1CD0] <= 0;
        weight_mem[16'h1CD1] <= 0;
        weight_mem[16'h1CD2] <= 0;
        weight_mem[16'h1CD3] <= 0;
        weight_mem[16'h1CD4] <= 0;
        weight_mem[16'h1CD5] <= 0;
        weight_mem[16'h1CD6] <= 0;
        weight_mem[16'h1CD7] <= 0;
        weight_mem[16'h1CD8] <= 0;
        weight_mem[16'h1CD9] <= 0;
        weight_mem[16'h1CDA] <= 0;
        weight_mem[16'h1CDB] <= 0;
        weight_mem[16'h1CDC] <= 0;
        weight_mem[16'h1CDD] <= 0;
        weight_mem[16'h1CDE] <= 0;
        weight_mem[16'h1CDF] <= 0;
        weight_mem[16'h1CE0] <= 0;
        weight_mem[16'h1CE1] <= 0;
        weight_mem[16'h1CE2] <= 0;
        weight_mem[16'h1CE3] <= 0;
        weight_mem[16'h1CE4] <= 0;
        weight_mem[16'h1CE5] <= 0;
        weight_mem[16'h1CE6] <= 0;
        weight_mem[16'h1CE7] <= 0;
        weight_mem[16'h1CE8] <= 0;
        weight_mem[16'h1CE9] <= 0;
        weight_mem[16'h1CEA] <= 0;
        weight_mem[16'h1CEB] <= 0;
        weight_mem[16'h1CEC] <= 0;
        weight_mem[16'h1CED] <= 0;
        weight_mem[16'h1CEE] <= 0;
        weight_mem[16'h1CEF] <= 0;
        weight_mem[16'h1CF0] <= 0;
        weight_mem[16'h1CF1] <= 0;
        weight_mem[16'h1CF2] <= 0;
        weight_mem[16'h1CF3] <= 0;
        weight_mem[16'h1CF4] <= 0;
        weight_mem[16'h1CF5] <= 0;
        weight_mem[16'h1CF6] <= 0;
        weight_mem[16'h1CF7] <= 0;
        weight_mem[16'h1CF8] <= 0;
        weight_mem[16'h1CF9] <= 0;
        weight_mem[16'h1CFA] <= 0;
        weight_mem[16'h1CFB] <= 0;
        weight_mem[16'h1CFC] <= 0;
        weight_mem[16'h1CFD] <= 0;
        weight_mem[16'h1CFE] <= 0;
        weight_mem[16'h1CFF] <= 0;
        weight_mem[16'h1D00] <= 0;
        weight_mem[16'h1D01] <= 0;
        weight_mem[16'h1D02] <= 0;
        weight_mem[16'h1D03] <= 0;
        weight_mem[16'h1D04] <= 0;
        weight_mem[16'h1D05] <= 0;
        weight_mem[16'h1D06] <= 0;
        weight_mem[16'h1D07] <= 0;
        weight_mem[16'h1D08] <= 0;
        weight_mem[16'h1D09] <= 0;
        weight_mem[16'h1D0A] <= 0;
        weight_mem[16'h1D0B] <= 0;
        weight_mem[16'h1D0C] <= 0;
        weight_mem[16'h1D0D] <= 0;
        weight_mem[16'h1D0E] <= 0;
        weight_mem[16'h1D0F] <= 0;
        weight_mem[16'h1D10] <= 0;
        weight_mem[16'h1D11] <= 0;
        weight_mem[16'h1D12] <= 0;
        weight_mem[16'h1D13] <= 0;
        weight_mem[16'h1D14] <= 0;
        weight_mem[16'h1D15] <= 0;
        weight_mem[16'h1D16] <= 0;
        weight_mem[16'h1D17] <= 0;
        weight_mem[16'h1D18] <= 0;
        weight_mem[16'h1D19] <= 0;
        weight_mem[16'h1D1A] <= 0;
        weight_mem[16'h1D1B] <= 0;
        weight_mem[16'h1D1C] <= 0;
        weight_mem[16'h1D1D] <= 0;
        weight_mem[16'h1D1E] <= 0;
        weight_mem[16'h1D1F] <= 0;
        weight_mem[16'h1D20] <= 0;
        weight_mem[16'h1D21] <= 0;
        weight_mem[16'h1D22] <= 0;
        weight_mem[16'h1D23] <= 0;
        weight_mem[16'h1D24] <= 0;
        weight_mem[16'h1D25] <= 0;
        weight_mem[16'h1D26] <= 0;
        weight_mem[16'h1D27] <= 0;
        weight_mem[16'h1D28] <= 0;
        weight_mem[16'h1D29] <= 0;
        weight_mem[16'h1D2A] <= 0;
        weight_mem[16'h1D2B] <= 0;
        weight_mem[16'h1D2C] <= 0;
        weight_mem[16'h1D2D] <= 0;
        weight_mem[16'h1D2E] <= 0;
        weight_mem[16'h1D2F] <= 0;
        weight_mem[16'h1D30] <= 0;
        weight_mem[16'h1D31] <= 0;
        weight_mem[16'h1D32] <= 0;
        weight_mem[16'h1D33] <= 0;
        weight_mem[16'h1D34] <= 0;
        weight_mem[16'h1D35] <= 0;
        weight_mem[16'h1D36] <= 0;
        weight_mem[16'h1D37] <= 0;
        weight_mem[16'h1D38] <= 0;
        weight_mem[16'h1D39] <= 0;
        weight_mem[16'h1D3A] <= 0;
        weight_mem[16'h1D3B] <= 0;
        weight_mem[16'h1D3C] <= 0;
        weight_mem[16'h1D3D] <= 0;
        weight_mem[16'h1D3E] <= 0;
        weight_mem[16'h1D3F] <= 0;
        weight_mem[16'h1D40] <= 0;
        weight_mem[16'h1D41] <= 0;
        weight_mem[16'h1D42] <= 0;
        weight_mem[16'h1D43] <= 0;
        weight_mem[16'h1D44] <= 0;
        weight_mem[16'h1D45] <= 0;
        weight_mem[16'h1D46] <= 0;
        weight_mem[16'h1D47] <= 0;
        weight_mem[16'h1D48] <= 0;
        weight_mem[16'h1D49] <= 0;
        weight_mem[16'h1D4A] <= 0;
        weight_mem[16'h1D4B] <= 0;
        weight_mem[16'h1D4C] <= 0;
        weight_mem[16'h1D4D] <= 0;
        weight_mem[16'h1D4E] <= 0;
        weight_mem[16'h1D4F] <= 0;
        weight_mem[16'h1D50] <= 0;
        weight_mem[16'h1D51] <= 0;
        weight_mem[16'h1D52] <= 0;
        weight_mem[16'h1D53] <= 0;
        weight_mem[16'h1D54] <= 0;
        weight_mem[16'h1D55] <= 0;
        weight_mem[16'h1D56] <= 0;
        weight_mem[16'h1D57] <= 0;
        weight_mem[16'h1D58] <= 0;
        weight_mem[16'h1D59] <= 0;
        weight_mem[16'h1D5A] <= 0;
        weight_mem[16'h1D5B] <= 0;
        weight_mem[16'h1D5C] <= 0;
        weight_mem[16'h1D5D] <= 0;
        weight_mem[16'h1D5E] <= 0;
        weight_mem[16'h1D5F] <= 0;
        weight_mem[16'h1D60] <= 0;
        weight_mem[16'h1D61] <= 0;
        weight_mem[16'h1D62] <= 0;
        weight_mem[16'h1D63] <= 0;
        weight_mem[16'h1D64] <= 0;
        weight_mem[16'h1D65] <= 0;
        weight_mem[16'h1D66] <= 0;
        weight_mem[16'h1D67] <= 0;
        weight_mem[16'h1D68] <= 0;
        weight_mem[16'h1D69] <= 0;
        weight_mem[16'h1D6A] <= 0;
        weight_mem[16'h1D6B] <= 0;
        weight_mem[16'h1D6C] <= 0;
        weight_mem[16'h1D6D] <= 0;
        weight_mem[16'h1D6E] <= 0;
        weight_mem[16'h1D6F] <= 0;
        weight_mem[16'h1D70] <= 0;
        weight_mem[16'h1D71] <= 0;
        weight_mem[16'h1D72] <= 0;
        weight_mem[16'h1D73] <= 0;
        weight_mem[16'h1D74] <= 0;
        weight_mem[16'h1D75] <= 0;
        weight_mem[16'h1D76] <= 0;
        weight_mem[16'h1D77] <= 0;
        weight_mem[16'h1D78] <= 0;
        weight_mem[16'h1D79] <= 0;
        weight_mem[16'h1D7A] <= 0;
        weight_mem[16'h1D7B] <= 0;
        weight_mem[16'h1D7C] <= 0;
        weight_mem[16'h1D7D] <= 0;
        weight_mem[16'h1D7E] <= 0;
        weight_mem[16'h1D7F] <= 0;
        weight_mem[16'h1D80] <= 0;
        weight_mem[16'h1D81] <= 0;
        weight_mem[16'h1D82] <= 0;
        weight_mem[16'h1D83] <= 0;
        weight_mem[16'h1D84] <= 0;
        weight_mem[16'h1D85] <= 0;
        weight_mem[16'h1D86] <= 0;
        weight_mem[16'h1D87] <= 0;
        weight_mem[16'h1D88] <= 0;
        weight_mem[16'h1D89] <= 0;
        weight_mem[16'h1D8A] <= 0;
        weight_mem[16'h1D8B] <= 0;
        weight_mem[16'h1D8C] <= 0;
        weight_mem[16'h1D8D] <= 0;
        weight_mem[16'h1D8E] <= 0;
        weight_mem[16'h1D8F] <= 0;
        weight_mem[16'h1D90] <= 0;
        weight_mem[16'h1D91] <= 0;
        weight_mem[16'h1D92] <= 0;
        weight_mem[16'h1D93] <= 0;
        weight_mem[16'h1D94] <= 0;
        weight_mem[16'h1D95] <= 0;
        weight_mem[16'h1D96] <= 0;
        weight_mem[16'h1D97] <= 0;
        weight_mem[16'h1D98] <= 0;
        weight_mem[16'h1D99] <= 0;
        weight_mem[16'h1D9A] <= 0;
        weight_mem[16'h1D9B] <= 0;
        weight_mem[16'h1D9C] <= 0;
        weight_mem[16'h1D9D] <= 0;
        weight_mem[16'h1D9E] <= 0;
        weight_mem[16'h1D9F] <= 0;
        weight_mem[16'h1DA0] <= 0;
        weight_mem[16'h1DA1] <= 0;
        weight_mem[16'h1DA2] <= 0;
        weight_mem[16'h1DA3] <= 0;
        weight_mem[16'h1DA4] <= 0;
        weight_mem[16'h1DA5] <= 0;
        weight_mem[16'h1DA6] <= 0;
        weight_mem[16'h1DA7] <= 0;
        weight_mem[16'h1DA8] <= 0;
        weight_mem[16'h1DA9] <= 0;
        weight_mem[16'h1DAA] <= 0;
        weight_mem[16'h1DAB] <= 0;
        weight_mem[16'h1DAC] <= 0;
        weight_mem[16'h1DAD] <= 0;
        weight_mem[16'h1DAE] <= 0;
        weight_mem[16'h1DAF] <= 0;

        // layer 1 neuron 15
        weight_mem[16'h1E00] <= 0;
        weight_mem[16'h1E01] <= 0;
        weight_mem[16'h1E02] <= 0;
        weight_mem[16'h1E03] <= 0;
        weight_mem[16'h1E04] <= 0;
        weight_mem[16'h1E05] <= 0;
        weight_mem[16'h1E06] <= 0;
        weight_mem[16'h1E07] <= 0;
        weight_mem[16'h1E08] <= 0;
        weight_mem[16'h1E09] <= 0;
        weight_mem[16'h1E0A] <= 0;
        weight_mem[16'h1E0B] <= 0;
        weight_mem[16'h1E0C] <= 0;
        weight_mem[16'h1E0D] <= 0;
        weight_mem[16'h1E0E] <= 0;
        weight_mem[16'h1E0F] <= 0;
        weight_mem[16'h1E10] <= 0;
        weight_mem[16'h1E11] <= 0;
        weight_mem[16'h1E12] <= 0;
        weight_mem[16'h1E13] <= 0;
        weight_mem[16'h1E14] <= 0;
        weight_mem[16'h1E15] <= 0;
        weight_mem[16'h1E16] <= 0;
        weight_mem[16'h1E17] <= 0;
        weight_mem[16'h1E18] <= 0;
        weight_mem[16'h1E19] <= 0;
        weight_mem[16'h1E1A] <= 0;
        weight_mem[16'h1E1B] <= 0;
        weight_mem[16'h1E1C] <= 0;
        weight_mem[16'h1E1D] <= 0;
        weight_mem[16'h1E1E] <= 0;
        weight_mem[16'h1E1F] <= 0;
        weight_mem[16'h1E20] <= 0;
        weight_mem[16'h1E21] <= 0;
        weight_mem[16'h1E22] <= 0;
        weight_mem[16'h1E23] <= 0;
        weight_mem[16'h1E24] <= 0;
        weight_mem[16'h1E25] <= 0;
        weight_mem[16'h1E26] <= 0;
        weight_mem[16'h1E27] <= 0;
        weight_mem[16'h1E28] <= 0;
        weight_mem[16'h1E29] <= 0;
        weight_mem[16'h1E2A] <= 0;
        weight_mem[16'h1E2B] <= 0;
        weight_mem[16'h1E2C] <= 0;
        weight_mem[16'h1E2D] <= 0;
        weight_mem[16'h1E2E] <= 0;
        weight_mem[16'h1E2F] <= 0;
        weight_mem[16'h1E30] <= 0;
        weight_mem[16'h1E31] <= 0;
        weight_mem[16'h1E32] <= 0;
        weight_mem[16'h1E33] <= 0;
        weight_mem[16'h1E34] <= 0;
        weight_mem[16'h1E35] <= 0;
        weight_mem[16'h1E36] <= 0;
        weight_mem[16'h1E37] <= 0;
        weight_mem[16'h1E38] <= 0;
        weight_mem[16'h1E39] <= 0;
        weight_mem[16'h1E3A] <= 0;
        weight_mem[16'h1E3B] <= 0;
        weight_mem[16'h1E3C] <= 0;
        weight_mem[16'h1E3D] <= 0;
        weight_mem[16'h1E3E] <= 0;
        weight_mem[16'h1E3F] <= 0;
        weight_mem[16'h1E40] <= 0;
        weight_mem[16'h1E41] <= 0;
        weight_mem[16'h1E42] <= 0;
        weight_mem[16'h1E43] <= 0;
        weight_mem[16'h1E44] <= 0;
        weight_mem[16'h1E45] <= 0;
        weight_mem[16'h1E46] <= 0;
        weight_mem[16'h1E47] <= 0;
        weight_mem[16'h1E48] <= 0;
        weight_mem[16'h1E49] <= 0;
        weight_mem[16'h1E4A] <= 0;
        weight_mem[16'h1E4B] <= 0;
        weight_mem[16'h1E4C] <= 0;
        weight_mem[16'h1E4D] <= 0;
        weight_mem[16'h1E4E] <= 0;
        weight_mem[16'h1E4F] <= 0;
        weight_mem[16'h1E50] <= 0;
        weight_mem[16'h1E51] <= 0;
        weight_mem[16'h1E52] <= 0;
        weight_mem[16'h1E53] <= 0;
        weight_mem[16'h1E54] <= 0;
        weight_mem[16'h1E55] <= 0;
        weight_mem[16'h1E56] <= 0;
        weight_mem[16'h1E57] <= 0;
        weight_mem[16'h1E58] <= 0;
        weight_mem[16'h1E59] <= 0;
        weight_mem[16'h1E5A] <= 0;
        weight_mem[16'h1E5B] <= 0;
        weight_mem[16'h1E5C] <= 0;
        weight_mem[16'h1E5D] <= 0;
        weight_mem[16'h1E5E] <= 0;
        weight_mem[16'h1E5F] <= 0;
        weight_mem[16'h1E60] <= 0;
        weight_mem[16'h1E61] <= 0;
        weight_mem[16'h1E62] <= 0;
        weight_mem[16'h1E63] <= 0;
        weight_mem[16'h1E64] <= 0;
        weight_mem[16'h1E65] <= 0;
        weight_mem[16'h1E66] <= 0;
        weight_mem[16'h1E67] <= 0;
        weight_mem[16'h1E68] <= 0;
        weight_mem[16'h1E69] <= 0;
        weight_mem[16'h1E6A] <= 0;
        weight_mem[16'h1E6B] <= 0;
        weight_mem[16'h1E6C] <= 0;
        weight_mem[16'h1E6D] <= 0;
        weight_mem[16'h1E6E] <= 0;
        weight_mem[16'h1E6F] <= 0;
        weight_mem[16'h1E70] <= 0;
        weight_mem[16'h1E71] <= 0;
        weight_mem[16'h1E72] <= 0;
        weight_mem[16'h1E73] <= 0;
        weight_mem[16'h1E74] <= 0;
        weight_mem[16'h1E75] <= 0;
        weight_mem[16'h1E76] <= 0;
        weight_mem[16'h1E77] <= 0;
        weight_mem[16'h1E78] <= 0;
        weight_mem[16'h1E79] <= 0;
        weight_mem[16'h1E7A] <= 0;
        weight_mem[16'h1E7B] <= 0;
        weight_mem[16'h1E7C] <= 0;
        weight_mem[16'h1E7D] <= 0;
        weight_mem[16'h1E7E] <= 0;
        weight_mem[16'h1E7F] <= 0;
        weight_mem[16'h1E80] <= 0;
        weight_mem[16'h1E81] <= 0;
        weight_mem[16'h1E82] <= 0;
        weight_mem[16'h1E83] <= 0;
        weight_mem[16'h1E84] <= 0;
        weight_mem[16'h1E85] <= 0;
        weight_mem[16'h1E86] <= 0;
        weight_mem[16'h1E87] <= 0;
        weight_mem[16'h1E88] <= 0;
        weight_mem[16'h1E89] <= 0;
        weight_mem[16'h1E8A] <= 0;
        weight_mem[16'h1E8B] <= 0;
        weight_mem[16'h1E8C] <= 0;
        weight_mem[16'h1E8D] <= 0;
        weight_mem[16'h1E8E] <= 0;
        weight_mem[16'h1E8F] <= 0;
        weight_mem[16'h1E90] <= 0;
        weight_mem[16'h1E91] <= 0;
        weight_mem[16'h1E92] <= 0;
        weight_mem[16'h1E93] <= 0;
        weight_mem[16'h1E94] <= 0;
        weight_mem[16'h1E95] <= 0;
        weight_mem[16'h1E96] <= 0;
        weight_mem[16'h1E97] <= 0;
        weight_mem[16'h1E98] <= 0;
        weight_mem[16'h1E99] <= 0;
        weight_mem[16'h1E9A] <= 0;
        weight_mem[16'h1E9B] <= 0;
        weight_mem[16'h1E9C] <= 0;
        weight_mem[16'h1E9D] <= 0;
        weight_mem[16'h1E9E] <= 0;
        weight_mem[16'h1E9F] <= 0;
        weight_mem[16'h1EA0] <= 0;
        weight_mem[16'h1EA1] <= 0;
        weight_mem[16'h1EA2] <= 0;
        weight_mem[16'h1EA3] <= 0;
        weight_mem[16'h1EA4] <= 0;
        weight_mem[16'h1EA5] <= 0;
        weight_mem[16'h1EA6] <= 0;
        weight_mem[16'h1EA7] <= 0;
        weight_mem[16'h1EA8] <= 0;
        weight_mem[16'h1EA9] <= 0;
        weight_mem[16'h1EAA] <= 0;
        weight_mem[16'h1EAB] <= 0;
        weight_mem[16'h1EAC] <= 0;
        weight_mem[16'h1EAD] <= 0;
        weight_mem[16'h1EAE] <= 0;
        weight_mem[16'h1EAF] <= 0;
        weight_mem[16'h1EB0] <= 0;
        weight_mem[16'h1EB1] <= 0;
        weight_mem[16'h1EB2] <= 0;
        weight_mem[16'h1EB3] <= 0;
        weight_mem[16'h1EB4] <= 0;
        weight_mem[16'h1EB5] <= 0;
        weight_mem[16'h1EB6] <= 0;
        weight_mem[16'h1EB7] <= 0;
        weight_mem[16'h1EB8] <= 0;
        weight_mem[16'h1EB9] <= 0;
        weight_mem[16'h1EBA] <= 0;
        weight_mem[16'h1EBB] <= 0;
        weight_mem[16'h1EBC] <= 0;
        weight_mem[16'h1EBD] <= 0;
        weight_mem[16'h1EBE] <= 0;
        weight_mem[16'h1EBF] <= 0;
        weight_mem[16'h1EC0] <= 0;
        weight_mem[16'h1EC1] <= 0;
        weight_mem[16'h1EC2] <= 0;
        weight_mem[16'h1EC3] <= 0;
        weight_mem[16'h1EC4] <= 0;
        weight_mem[16'h1EC5] <= 0;
        weight_mem[16'h1EC6] <= 0;
        weight_mem[16'h1EC7] <= 0;
        weight_mem[16'h1EC8] <= 0;
        weight_mem[16'h1EC9] <= 0;
        weight_mem[16'h1ECA] <= 0;
        weight_mem[16'h1ECB] <= 0;
        weight_mem[16'h1ECC] <= 0;
        weight_mem[16'h1ECD] <= 0;
        weight_mem[16'h1ECE] <= 0;
        weight_mem[16'h1ECF] <= 0;
        weight_mem[16'h1ED0] <= 0;
        weight_mem[16'h1ED1] <= 0;
        weight_mem[16'h1ED2] <= 0;
        weight_mem[16'h1ED3] <= 0;
        weight_mem[16'h1ED4] <= 0;
        weight_mem[16'h1ED5] <= 0;
        weight_mem[16'h1ED6] <= 0;
        weight_mem[16'h1ED7] <= 0;
        weight_mem[16'h1ED8] <= 0;
        weight_mem[16'h1ED9] <= 0;
        weight_mem[16'h1EDA] <= 0;
        weight_mem[16'h1EDB] <= 0;
        weight_mem[16'h1EDC] <= 0;
        weight_mem[16'h1EDD] <= 0;
        weight_mem[16'h1EDE] <= 0;
        weight_mem[16'h1EDF] <= 0;
        weight_mem[16'h1EE0] <= 0;
        weight_mem[16'h1EE1] <= 0;
        weight_mem[16'h1EE2] <= 0;
        weight_mem[16'h1EE3] <= 0;
        weight_mem[16'h1EE4] <= 0;
        weight_mem[16'h1EE5] <= 0;
        weight_mem[16'h1EE6] <= 0;
        weight_mem[16'h1EE7] <= 0;
        weight_mem[16'h1EE8] <= 0;
        weight_mem[16'h1EE9] <= 0;
        weight_mem[16'h1EEA] <= 0;
        weight_mem[16'h1EEB] <= 0;
        weight_mem[16'h1EEC] <= 0;
        weight_mem[16'h1EED] <= 0;
        weight_mem[16'h1EEE] <= 0;
        weight_mem[16'h1EEF] <= 0;
        weight_mem[16'h1EF0] <= 0;
        weight_mem[16'h1EF1] <= 0;
        weight_mem[16'h1EF2] <= 0;
        weight_mem[16'h1EF3] <= 0;
        weight_mem[16'h1EF4] <= 0;
        weight_mem[16'h1EF5] <= 0;
        weight_mem[16'h1EF6] <= 0;
        weight_mem[16'h1EF7] <= 0;
        weight_mem[16'h1EF8] <= 0;
        weight_mem[16'h1EF9] <= 0;
        weight_mem[16'h1EFA] <= 0;
        weight_mem[16'h1EFB] <= 0;
        weight_mem[16'h1EFC] <= 0;
        weight_mem[16'h1EFD] <= 0;
        weight_mem[16'h1EFE] <= 0;
        weight_mem[16'h1EFF] <= 0;
        weight_mem[16'h1F00] <= 0;
        weight_mem[16'h1F01] <= 0;
        weight_mem[16'h1F02] <= 0;
        weight_mem[16'h1F03] <= 0;
        weight_mem[16'h1F04] <= 0;
        weight_mem[16'h1F05] <= 0;
        weight_mem[16'h1F06] <= 0;
        weight_mem[16'h1F07] <= 0;
        weight_mem[16'h1F08] <= 0;
        weight_mem[16'h1F09] <= 0;
        weight_mem[16'h1F0A] <= 0;
        weight_mem[16'h1F0B] <= 0;
        weight_mem[16'h1F0C] <= 0;
        weight_mem[16'h1F0D] <= 0;
        weight_mem[16'h1F0E] <= 0;
        weight_mem[16'h1F0F] <= 0;
        weight_mem[16'h1F10] <= 0;
        weight_mem[16'h1F11] <= 0;
        weight_mem[16'h1F12] <= 0;
        weight_mem[16'h1F13] <= 0;
        weight_mem[16'h1F14] <= 0;
        weight_mem[16'h1F15] <= 0;
        weight_mem[16'h1F16] <= 0;
        weight_mem[16'h1F17] <= 0;
        weight_mem[16'h1F18] <= 0;
        weight_mem[16'h1F19] <= 0;
        weight_mem[16'h1F1A] <= 0;
        weight_mem[16'h1F1B] <= 0;
        weight_mem[16'h1F1C] <= 0;
        weight_mem[16'h1F1D] <= 0;
        weight_mem[16'h1F1E] <= 0;
        weight_mem[16'h1F1F] <= 0;
        weight_mem[16'h1F20] <= 0;
        weight_mem[16'h1F21] <= 0;
        weight_mem[16'h1F22] <= 0;
        weight_mem[16'h1F23] <= 0;
        weight_mem[16'h1F24] <= 0;
        weight_mem[16'h1F25] <= 0;
        weight_mem[16'h1F26] <= 0;
        weight_mem[16'h1F27] <= 0;
        weight_mem[16'h1F28] <= 0;
        weight_mem[16'h1F29] <= 0;
        weight_mem[16'h1F2A] <= 0;
        weight_mem[16'h1F2B] <= 0;
        weight_mem[16'h1F2C] <= 0;
        weight_mem[16'h1F2D] <= 0;
        weight_mem[16'h1F2E] <= 0;
        weight_mem[16'h1F2F] <= 0;
        weight_mem[16'h1F30] <= 0;
        weight_mem[16'h1F31] <= 0;
        weight_mem[16'h1F32] <= 0;
        weight_mem[16'h1F33] <= 0;
        weight_mem[16'h1F34] <= 0;
        weight_mem[16'h1F35] <= 0;
        weight_mem[16'h1F36] <= 0;
        weight_mem[16'h1F37] <= 0;
        weight_mem[16'h1F38] <= 0;
        weight_mem[16'h1F39] <= 0;
        weight_mem[16'h1F3A] <= 0;
        weight_mem[16'h1F3B] <= 0;
        weight_mem[16'h1F3C] <= 0;
        weight_mem[16'h1F3D] <= 0;
        weight_mem[16'h1F3E] <= 0;
        weight_mem[16'h1F3F] <= 0;
        weight_mem[16'h1F40] <= 0;
        weight_mem[16'h1F41] <= 0;
        weight_mem[16'h1F42] <= 0;
        weight_mem[16'h1F43] <= 0;
        weight_mem[16'h1F44] <= 0;
        weight_mem[16'h1F45] <= 0;
        weight_mem[16'h1F46] <= 0;
        weight_mem[16'h1F47] <= 0;
        weight_mem[16'h1F48] <= 0;
        weight_mem[16'h1F49] <= 0;
        weight_mem[16'h1F4A] <= 0;
        weight_mem[16'h1F4B] <= 0;
        weight_mem[16'h1F4C] <= 0;
        weight_mem[16'h1F4D] <= 0;
        weight_mem[16'h1F4E] <= 0;
        weight_mem[16'h1F4F] <= 0;
        weight_mem[16'h1F50] <= 0;
        weight_mem[16'h1F51] <= 0;
        weight_mem[16'h1F52] <= 0;
        weight_mem[16'h1F53] <= 0;
        weight_mem[16'h1F54] <= 0;
        weight_mem[16'h1F55] <= 0;
        weight_mem[16'h1F56] <= 0;
        weight_mem[16'h1F57] <= 0;
        weight_mem[16'h1F58] <= 0;
        weight_mem[16'h1F59] <= 0;
        weight_mem[16'h1F5A] <= 0;
        weight_mem[16'h1F5B] <= 0;
        weight_mem[16'h1F5C] <= 0;
        weight_mem[16'h1F5D] <= 0;
        weight_mem[16'h1F5E] <= 0;
        weight_mem[16'h1F5F] <= 0;
        weight_mem[16'h1F60] <= 0;
        weight_mem[16'h1F61] <= 0;
        weight_mem[16'h1F62] <= 0;
        weight_mem[16'h1F63] <= 0;
        weight_mem[16'h1F64] <= 0;
        weight_mem[16'h1F65] <= 0;
        weight_mem[16'h1F66] <= 0;
        weight_mem[16'h1F67] <= 0;
        weight_mem[16'h1F68] <= 0;
        weight_mem[16'h1F69] <= 0;
        weight_mem[16'h1F6A] <= 0;
        weight_mem[16'h1F6B] <= 0;
        weight_mem[16'h1F6C] <= 0;
        weight_mem[16'h1F6D] <= 0;
        weight_mem[16'h1F6E] <= 0;
        weight_mem[16'h1F6F] <= 0;
        weight_mem[16'h1F70] <= 0;
        weight_mem[16'h1F71] <= 0;
        weight_mem[16'h1F72] <= 0;
        weight_mem[16'h1F73] <= 0;
        weight_mem[16'h1F74] <= 0;
        weight_mem[16'h1F75] <= 0;
        weight_mem[16'h1F76] <= 0;
        weight_mem[16'h1F77] <= 0;
        weight_mem[16'h1F78] <= 0;
        weight_mem[16'h1F79] <= 0;
        weight_mem[16'h1F7A] <= 0;
        weight_mem[16'h1F7B] <= 0;
        weight_mem[16'h1F7C] <= 0;
        weight_mem[16'h1F7D] <= 0;
        weight_mem[16'h1F7E] <= 0;
        weight_mem[16'h1F7F] <= 0;
        weight_mem[16'h1F80] <= 0;
        weight_mem[16'h1F81] <= 0;
        weight_mem[16'h1F82] <= 0;
        weight_mem[16'h1F83] <= 0;
        weight_mem[16'h1F84] <= 0;
        weight_mem[16'h1F85] <= 0;
        weight_mem[16'h1F86] <= 0;
        weight_mem[16'h1F87] <= 0;
        weight_mem[16'h1F88] <= 0;
        weight_mem[16'h1F89] <= 0;
        weight_mem[16'h1F8A] <= 0;
        weight_mem[16'h1F8B] <= 0;
        weight_mem[16'h1F8C] <= 0;
        weight_mem[16'h1F8D] <= 0;
        weight_mem[16'h1F8E] <= 0;
        weight_mem[16'h1F8F] <= 0;
        weight_mem[16'h1F90] <= 0;
        weight_mem[16'h1F91] <= 0;
        weight_mem[16'h1F92] <= 0;
        weight_mem[16'h1F93] <= 0;
        weight_mem[16'h1F94] <= 0;
        weight_mem[16'h1F95] <= 0;
        weight_mem[16'h1F96] <= 0;
        weight_mem[16'h1F97] <= 0;
        weight_mem[16'h1F98] <= 0;
        weight_mem[16'h1F99] <= 0;
        weight_mem[16'h1F9A] <= 0;
        weight_mem[16'h1F9B] <= 0;
        weight_mem[16'h1F9C] <= 0;
        weight_mem[16'h1F9D] <= 0;
        weight_mem[16'h1F9E] <= 0;
        weight_mem[16'h1F9F] <= 0;
        weight_mem[16'h1FA0] <= 0;
        weight_mem[16'h1FA1] <= 0;
        weight_mem[16'h1FA2] <= 0;
        weight_mem[16'h1FA3] <= 0;
        weight_mem[16'h1FA4] <= 0;
        weight_mem[16'h1FA5] <= 0;
        weight_mem[16'h1FA6] <= 0;
        weight_mem[16'h1FA7] <= 0;
        weight_mem[16'h1FA8] <= 0;
        weight_mem[16'h1FA9] <= 0;
        weight_mem[16'h1FAA] <= 0;
        weight_mem[16'h1FAB] <= 0;
        weight_mem[16'h1FAC] <= 0;
        weight_mem[16'h1FAD] <= 0;
        weight_mem[16'h1FAE] <= 0;
        weight_mem[16'h1FAF] <= 0;

        // layer 1 neuron 16
        weight_mem[16'h2000] <= 0;
        weight_mem[16'h2001] <= 0;
        weight_mem[16'h2002] <= 0;
        weight_mem[16'h2003] <= 0;
        weight_mem[16'h2004] <= 0;
        weight_mem[16'h2005] <= 0;
        weight_mem[16'h2006] <= 0;
        weight_mem[16'h2007] <= 0;
        weight_mem[16'h2008] <= 0;
        weight_mem[16'h2009] <= 0;
        weight_mem[16'h200A] <= 0;
        weight_mem[16'h200B] <= 0;
        weight_mem[16'h200C] <= 0;
        weight_mem[16'h200D] <= 0;
        weight_mem[16'h200E] <= 0;
        weight_mem[16'h200F] <= 0;
        weight_mem[16'h2010] <= 0;
        weight_mem[16'h2011] <= 0;
        weight_mem[16'h2012] <= 0;
        weight_mem[16'h2013] <= 0;
        weight_mem[16'h2014] <= 0;
        weight_mem[16'h2015] <= 0;
        weight_mem[16'h2016] <= 0;
        weight_mem[16'h2017] <= 0;
        weight_mem[16'h2018] <= 0;
        weight_mem[16'h2019] <= 0;
        weight_mem[16'h201A] <= 0;
        weight_mem[16'h201B] <= 0;
        weight_mem[16'h201C] <= 0;
        weight_mem[16'h201D] <= 0;
        weight_mem[16'h201E] <= 0;
        weight_mem[16'h201F] <= 0;
        weight_mem[16'h2020] <= 0;
        weight_mem[16'h2021] <= 0;
        weight_mem[16'h2022] <= 0;
        weight_mem[16'h2023] <= 0;
        weight_mem[16'h2024] <= 0;
        weight_mem[16'h2025] <= 0;
        weight_mem[16'h2026] <= 0;
        weight_mem[16'h2027] <= 0;
        weight_mem[16'h2028] <= 0;
        weight_mem[16'h2029] <= 0;
        weight_mem[16'h202A] <= 0;
        weight_mem[16'h202B] <= 0;
        weight_mem[16'h202C] <= 0;
        weight_mem[16'h202D] <= 0;
        weight_mem[16'h202E] <= 0;
        weight_mem[16'h202F] <= 0;
        weight_mem[16'h2030] <= 0;
        weight_mem[16'h2031] <= 0;
        weight_mem[16'h2032] <= 0;
        weight_mem[16'h2033] <= 0;
        weight_mem[16'h2034] <= 0;
        weight_mem[16'h2035] <= 0;
        weight_mem[16'h2036] <= 0;
        weight_mem[16'h2037] <= 0;
        weight_mem[16'h2038] <= 0;
        weight_mem[16'h2039] <= 0;
        weight_mem[16'h203A] <= 0;
        weight_mem[16'h203B] <= 0;
        weight_mem[16'h203C] <= 0;
        weight_mem[16'h203D] <= 0;
        weight_mem[16'h203E] <= 0;
        weight_mem[16'h203F] <= 0;
        weight_mem[16'h2040] <= 0;
        weight_mem[16'h2041] <= 0;
        weight_mem[16'h2042] <= 0;
        weight_mem[16'h2043] <= 0;
        weight_mem[16'h2044] <= 0;
        weight_mem[16'h2045] <= 0;
        weight_mem[16'h2046] <= 0;
        weight_mem[16'h2047] <= 0;
        weight_mem[16'h2048] <= 0;
        weight_mem[16'h2049] <= 0;
        weight_mem[16'h204A] <= 0;
        weight_mem[16'h204B] <= 0;
        weight_mem[16'h204C] <= 0;
        weight_mem[16'h204D] <= 0;
        weight_mem[16'h204E] <= 0;
        weight_mem[16'h204F] <= 0;
        weight_mem[16'h2050] <= 0;
        weight_mem[16'h2051] <= 0;
        weight_mem[16'h2052] <= 0;
        weight_mem[16'h2053] <= 0;
        weight_mem[16'h2054] <= 0;
        weight_mem[16'h2055] <= 0;
        weight_mem[16'h2056] <= 0;
        weight_mem[16'h2057] <= 0;
        weight_mem[16'h2058] <= 0;
        weight_mem[16'h2059] <= 0;
        weight_mem[16'h205A] <= 0;
        weight_mem[16'h205B] <= 0;
        weight_mem[16'h205C] <= 0;
        weight_mem[16'h205D] <= 0;
        weight_mem[16'h205E] <= 0;
        weight_mem[16'h205F] <= 0;
        weight_mem[16'h2060] <= 0;
        weight_mem[16'h2061] <= 0;
        weight_mem[16'h2062] <= 0;
        weight_mem[16'h2063] <= 0;
        weight_mem[16'h2064] <= 0;
        weight_mem[16'h2065] <= 0;
        weight_mem[16'h2066] <= 0;
        weight_mem[16'h2067] <= 0;
        weight_mem[16'h2068] <= 0;
        weight_mem[16'h2069] <= 0;
        weight_mem[16'h206A] <= 0;
        weight_mem[16'h206B] <= 0;
        weight_mem[16'h206C] <= 0;
        weight_mem[16'h206D] <= 0;
        weight_mem[16'h206E] <= 0;
        weight_mem[16'h206F] <= 0;
        weight_mem[16'h2070] <= 0;
        weight_mem[16'h2071] <= 0;
        weight_mem[16'h2072] <= 0;
        weight_mem[16'h2073] <= 0;
        weight_mem[16'h2074] <= 0;
        weight_mem[16'h2075] <= 0;
        weight_mem[16'h2076] <= 0;
        weight_mem[16'h2077] <= 0;
        weight_mem[16'h2078] <= 0;
        weight_mem[16'h2079] <= 0;
        weight_mem[16'h207A] <= 0;
        weight_mem[16'h207B] <= 0;
        weight_mem[16'h207C] <= 0;
        weight_mem[16'h207D] <= 0;
        weight_mem[16'h207E] <= 0;
        weight_mem[16'h207F] <= 0;
        weight_mem[16'h2080] <= 0;
        weight_mem[16'h2081] <= 0;
        weight_mem[16'h2082] <= 0;
        weight_mem[16'h2083] <= 0;
        weight_mem[16'h2084] <= 0;
        weight_mem[16'h2085] <= 0;
        weight_mem[16'h2086] <= 0;
        weight_mem[16'h2087] <= 0;
        weight_mem[16'h2088] <= 0;
        weight_mem[16'h2089] <= 0;
        weight_mem[16'h208A] <= 0;
        weight_mem[16'h208B] <= 0;
        weight_mem[16'h208C] <= 0;
        weight_mem[16'h208D] <= 0;
        weight_mem[16'h208E] <= 0;
        weight_mem[16'h208F] <= 0;
        weight_mem[16'h2090] <= 0;
        weight_mem[16'h2091] <= 0;
        weight_mem[16'h2092] <= 0;
        weight_mem[16'h2093] <= 0;
        weight_mem[16'h2094] <= 0;
        weight_mem[16'h2095] <= 0;
        weight_mem[16'h2096] <= 0;
        weight_mem[16'h2097] <= 0;
        weight_mem[16'h2098] <= 0;
        weight_mem[16'h2099] <= 0;
        weight_mem[16'h209A] <= 0;
        weight_mem[16'h209B] <= 0;
        weight_mem[16'h209C] <= 0;
        weight_mem[16'h209D] <= 0;
        weight_mem[16'h209E] <= 0;
        weight_mem[16'h209F] <= 0;
        weight_mem[16'h20A0] <= 0;
        weight_mem[16'h20A1] <= 0;
        weight_mem[16'h20A2] <= 0;
        weight_mem[16'h20A3] <= 0;
        weight_mem[16'h20A4] <= 0;
        weight_mem[16'h20A5] <= 0;
        weight_mem[16'h20A6] <= 0;
        weight_mem[16'h20A7] <= 0;
        weight_mem[16'h20A8] <= 0;
        weight_mem[16'h20A9] <= 0;
        weight_mem[16'h20AA] <= 0;
        weight_mem[16'h20AB] <= 0;
        weight_mem[16'h20AC] <= 0;
        weight_mem[16'h20AD] <= 0;
        weight_mem[16'h20AE] <= 0;
        weight_mem[16'h20AF] <= 0;
        weight_mem[16'h20B0] <= 0;
        weight_mem[16'h20B1] <= 0;
        weight_mem[16'h20B2] <= 0;
        weight_mem[16'h20B3] <= 0;
        weight_mem[16'h20B4] <= 0;
        weight_mem[16'h20B5] <= 0;
        weight_mem[16'h20B6] <= 0;
        weight_mem[16'h20B7] <= 0;
        weight_mem[16'h20B8] <= 0;
        weight_mem[16'h20B9] <= 0;
        weight_mem[16'h20BA] <= 0;
        weight_mem[16'h20BB] <= 0;
        weight_mem[16'h20BC] <= 0;
        weight_mem[16'h20BD] <= 0;
        weight_mem[16'h20BE] <= 0;
        weight_mem[16'h20BF] <= 0;
        weight_mem[16'h20C0] <= 0;
        weight_mem[16'h20C1] <= 0;
        weight_mem[16'h20C2] <= 0;
        weight_mem[16'h20C3] <= 0;
        weight_mem[16'h20C4] <= 0;
        weight_mem[16'h20C5] <= 0;
        weight_mem[16'h20C6] <= 0;
        weight_mem[16'h20C7] <= 0;
        weight_mem[16'h20C8] <= 0;
        weight_mem[16'h20C9] <= 0;
        weight_mem[16'h20CA] <= 0;
        weight_mem[16'h20CB] <= 0;
        weight_mem[16'h20CC] <= 0;
        weight_mem[16'h20CD] <= 0;
        weight_mem[16'h20CE] <= 0;
        weight_mem[16'h20CF] <= 0;
        weight_mem[16'h20D0] <= 0;
        weight_mem[16'h20D1] <= 0;
        weight_mem[16'h20D2] <= 0;
        weight_mem[16'h20D3] <= 0;
        weight_mem[16'h20D4] <= 0;
        weight_mem[16'h20D5] <= 0;
        weight_mem[16'h20D6] <= 0;
        weight_mem[16'h20D7] <= 0;
        weight_mem[16'h20D8] <= 0;
        weight_mem[16'h20D9] <= 0;
        weight_mem[16'h20DA] <= 0;
        weight_mem[16'h20DB] <= 0;
        weight_mem[16'h20DC] <= 0;
        weight_mem[16'h20DD] <= 0;
        weight_mem[16'h20DE] <= 0;
        weight_mem[16'h20DF] <= 0;
        weight_mem[16'h20E0] <= 0;
        weight_mem[16'h20E1] <= 0;
        weight_mem[16'h20E2] <= 0;
        weight_mem[16'h20E3] <= 0;
        weight_mem[16'h20E4] <= 0;
        weight_mem[16'h20E5] <= 0;
        weight_mem[16'h20E6] <= 0;
        weight_mem[16'h20E7] <= 0;
        weight_mem[16'h20E8] <= 0;
        weight_mem[16'h20E9] <= 0;
        weight_mem[16'h20EA] <= 0;
        weight_mem[16'h20EB] <= 0;
        weight_mem[16'h20EC] <= 0;
        weight_mem[16'h20ED] <= 0;
        weight_mem[16'h20EE] <= 0;
        weight_mem[16'h20EF] <= 0;
        weight_mem[16'h20F0] <= 0;
        weight_mem[16'h20F1] <= 0;
        weight_mem[16'h20F2] <= 0;
        weight_mem[16'h20F3] <= 0;
        weight_mem[16'h20F4] <= 0;
        weight_mem[16'h20F5] <= 0;
        weight_mem[16'h20F6] <= 0;
        weight_mem[16'h20F7] <= 0;
        weight_mem[16'h20F8] <= 0;
        weight_mem[16'h20F9] <= 0;
        weight_mem[16'h20FA] <= 0;
        weight_mem[16'h20FB] <= 0;
        weight_mem[16'h20FC] <= 0;
        weight_mem[16'h20FD] <= 0;
        weight_mem[16'h20FE] <= 0;
        weight_mem[16'h20FF] <= 0;
        weight_mem[16'h2100] <= 0;
        weight_mem[16'h2101] <= 0;
        weight_mem[16'h2102] <= 0;
        weight_mem[16'h2103] <= 0;
        weight_mem[16'h2104] <= 0;
        weight_mem[16'h2105] <= 0;
        weight_mem[16'h2106] <= 0;
        weight_mem[16'h2107] <= 0;
        weight_mem[16'h2108] <= 0;
        weight_mem[16'h2109] <= 0;
        weight_mem[16'h210A] <= 0;
        weight_mem[16'h210B] <= 0;
        weight_mem[16'h210C] <= 0;
        weight_mem[16'h210D] <= 0;
        weight_mem[16'h210E] <= 0;
        weight_mem[16'h210F] <= 0;
        weight_mem[16'h2110] <= 0;
        weight_mem[16'h2111] <= 0;
        weight_mem[16'h2112] <= 0;
        weight_mem[16'h2113] <= 0;
        weight_mem[16'h2114] <= 0;
        weight_mem[16'h2115] <= 0;
        weight_mem[16'h2116] <= 0;
        weight_mem[16'h2117] <= 0;
        weight_mem[16'h2118] <= 0;
        weight_mem[16'h2119] <= 0;
        weight_mem[16'h211A] <= 0;
        weight_mem[16'h211B] <= 0;
        weight_mem[16'h211C] <= 0;
        weight_mem[16'h211D] <= 0;
        weight_mem[16'h211E] <= 0;
        weight_mem[16'h211F] <= 0;
        weight_mem[16'h2120] <= 0;
        weight_mem[16'h2121] <= 0;
        weight_mem[16'h2122] <= 0;
        weight_mem[16'h2123] <= 0;
        weight_mem[16'h2124] <= 0;
        weight_mem[16'h2125] <= 0;
        weight_mem[16'h2126] <= 0;
        weight_mem[16'h2127] <= 0;
        weight_mem[16'h2128] <= 0;
        weight_mem[16'h2129] <= 0;
        weight_mem[16'h212A] <= 0;
        weight_mem[16'h212B] <= 0;
        weight_mem[16'h212C] <= 0;
        weight_mem[16'h212D] <= 0;
        weight_mem[16'h212E] <= 0;
        weight_mem[16'h212F] <= 0;
        weight_mem[16'h2130] <= 0;
        weight_mem[16'h2131] <= 0;
        weight_mem[16'h2132] <= 0;
        weight_mem[16'h2133] <= 0;
        weight_mem[16'h2134] <= 0;
        weight_mem[16'h2135] <= 0;
        weight_mem[16'h2136] <= 0;
        weight_mem[16'h2137] <= 0;
        weight_mem[16'h2138] <= 0;
        weight_mem[16'h2139] <= 0;
        weight_mem[16'h213A] <= 0;
        weight_mem[16'h213B] <= 0;
        weight_mem[16'h213C] <= 0;
        weight_mem[16'h213D] <= 0;
        weight_mem[16'h213E] <= 0;
        weight_mem[16'h213F] <= 0;
        weight_mem[16'h2140] <= 0;
        weight_mem[16'h2141] <= 0;
        weight_mem[16'h2142] <= 0;
        weight_mem[16'h2143] <= 0;
        weight_mem[16'h2144] <= 0;
        weight_mem[16'h2145] <= 0;
        weight_mem[16'h2146] <= 0;
        weight_mem[16'h2147] <= 0;
        weight_mem[16'h2148] <= 0;
        weight_mem[16'h2149] <= 0;
        weight_mem[16'h214A] <= 0;
        weight_mem[16'h214B] <= 0;
        weight_mem[16'h214C] <= 0;
        weight_mem[16'h214D] <= 0;
        weight_mem[16'h214E] <= 0;
        weight_mem[16'h214F] <= 0;
        weight_mem[16'h2150] <= 0;
        weight_mem[16'h2151] <= 0;
        weight_mem[16'h2152] <= 0;
        weight_mem[16'h2153] <= 0;
        weight_mem[16'h2154] <= 0;
        weight_mem[16'h2155] <= 0;
        weight_mem[16'h2156] <= 0;
        weight_mem[16'h2157] <= 0;
        weight_mem[16'h2158] <= 0;
        weight_mem[16'h2159] <= 0;
        weight_mem[16'h215A] <= 0;
        weight_mem[16'h215B] <= 0;
        weight_mem[16'h215C] <= 0;
        weight_mem[16'h215D] <= 0;
        weight_mem[16'h215E] <= 0;
        weight_mem[16'h215F] <= 0;
        weight_mem[16'h2160] <= 0;
        weight_mem[16'h2161] <= 0;
        weight_mem[16'h2162] <= 0;
        weight_mem[16'h2163] <= 0;
        weight_mem[16'h2164] <= 0;
        weight_mem[16'h2165] <= 0;
        weight_mem[16'h2166] <= 0;
        weight_mem[16'h2167] <= 0;
        weight_mem[16'h2168] <= 0;
        weight_mem[16'h2169] <= 0;
        weight_mem[16'h216A] <= 0;
        weight_mem[16'h216B] <= 0;
        weight_mem[16'h216C] <= 0;
        weight_mem[16'h216D] <= 0;
        weight_mem[16'h216E] <= 0;
        weight_mem[16'h216F] <= 0;
        weight_mem[16'h2170] <= 0;
        weight_mem[16'h2171] <= 0;
        weight_mem[16'h2172] <= 0;
        weight_mem[16'h2173] <= 0;
        weight_mem[16'h2174] <= 0;
        weight_mem[16'h2175] <= 0;
        weight_mem[16'h2176] <= 0;
        weight_mem[16'h2177] <= 0;
        weight_mem[16'h2178] <= 0;
        weight_mem[16'h2179] <= 0;
        weight_mem[16'h217A] <= 0;
        weight_mem[16'h217B] <= 0;
        weight_mem[16'h217C] <= 0;
        weight_mem[16'h217D] <= 0;
        weight_mem[16'h217E] <= 0;
        weight_mem[16'h217F] <= 0;
        weight_mem[16'h2180] <= 0;
        weight_mem[16'h2181] <= 0;
        weight_mem[16'h2182] <= 0;
        weight_mem[16'h2183] <= 0;
        weight_mem[16'h2184] <= 0;
        weight_mem[16'h2185] <= 0;
        weight_mem[16'h2186] <= 0;
        weight_mem[16'h2187] <= 0;
        weight_mem[16'h2188] <= 0;
        weight_mem[16'h2189] <= 0;
        weight_mem[16'h218A] <= 0;
        weight_mem[16'h218B] <= 0;
        weight_mem[16'h218C] <= 0;
        weight_mem[16'h218D] <= 0;
        weight_mem[16'h218E] <= 0;
        weight_mem[16'h218F] <= 0;
        weight_mem[16'h2190] <= 0;
        weight_mem[16'h2191] <= 0;
        weight_mem[16'h2192] <= 0;
        weight_mem[16'h2193] <= 0;
        weight_mem[16'h2194] <= 0;
        weight_mem[16'h2195] <= 0;
        weight_mem[16'h2196] <= 0;
        weight_mem[16'h2197] <= 0;
        weight_mem[16'h2198] <= 0;
        weight_mem[16'h2199] <= 0;
        weight_mem[16'h219A] <= 0;
        weight_mem[16'h219B] <= 0;
        weight_mem[16'h219C] <= 0;
        weight_mem[16'h219D] <= 0;
        weight_mem[16'h219E] <= 0;
        weight_mem[16'h219F] <= 0;
        weight_mem[16'h21A0] <= 0;
        weight_mem[16'h21A1] <= 0;
        weight_mem[16'h21A2] <= 0;
        weight_mem[16'h21A3] <= 0;
        weight_mem[16'h21A4] <= 0;
        weight_mem[16'h21A5] <= 0;
        weight_mem[16'h21A6] <= 0;
        weight_mem[16'h21A7] <= 0;
        weight_mem[16'h21A8] <= 0;
        weight_mem[16'h21A9] <= 0;
        weight_mem[16'h21AA] <= 0;
        weight_mem[16'h21AB] <= 0;
        weight_mem[16'h21AC] <= 0;
        weight_mem[16'h21AD] <= 0;
        weight_mem[16'h21AE] <= 0;
        weight_mem[16'h21AF] <= 0;

        // layer 1 neuron 17
        weight_mem[16'h2200] <= 0;
        weight_mem[16'h2201] <= 0;
        weight_mem[16'h2202] <= 0;
        weight_mem[16'h2203] <= 0;
        weight_mem[16'h2204] <= 0;
        weight_mem[16'h2205] <= 0;
        weight_mem[16'h2206] <= 0;
        weight_mem[16'h2207] <= 0;
        weight_mem[16'h2208] <= 0;
        weight_mem[16'h2209] <= 0;
        weight_mem[16'h220A] <= 0;
        weight_mem[16'h220B] <= 0;
        weight_mem[16'h220C] <= 0;
        weight_mem[16'h220D] <= 0;
        weight_mem[16'h220E] <= 0;
        weight_mem[16'h220F] <= 0;
        weight_mem[16'h2210] <= 0;
        weight_mem[16'h2211] <= 0;
        weight_mem[16'h2212] <= 0;
        weight_mem[16'h2213] <= 0;
        weight_mem[16'h2214] <= 0;
        weight_mem[16'h2215] <= 0;
        weight_mem[16'h2216] <= 0;
        weight_mem[16'h2217] <= 0;
        weight_mem[16'h2218] <= 0;
        weight_mem[16'h2219] <= 0;
        weight_mem[16'h221A] <= 0;
        weight_mem[16'h221B] <= 0;
        weight_mem[16'h221C] <= 0;
        weight_mem[16'h221D] <= 0;
        weight_mem[16'h221E] <= 0;
        weight_mem[16'h221F] <= 0;
        weight_mem[16'h2220] <= 0;
        weight_mem[16'h2221] <= 0;
        weight_mem[16'h2222] <= 0;
        weight_mem[16'h2223] <= 0;
        weight_mem[16'h2224] <= 0;
        weight_mem[16'h2225] <= 0;
        weight_mem[16'h2226] <= 0;
        weight_mem[16'h2227] <= 0;
        weight_mem[16'h2228] <= 0;
        weight_mem[16'h2229] <= 0;
        weight_mem[16'h222A] <= 0;
        weight_mem[16'h222B] <= 0;
        weight_mem[16'h222C] <= 0;
        weight_mem[16'h222D] <= 0;
        weight_mem[16'h222E] <= 0;
        weight_mem[16'h222F] <= 0;
        weight_mem[16'h2230] <= 0;
        weight_mem[16'h2231] <= 0;
        weight_mem[16'h2232] <= 0;
        weight_mem[16'h2233] <= 0;
        weight_mem[16'h2234] <= 0;
        weight_mem[16'h2235] <= 0;
        weight_mem[16'h2236] <= 0;
        weight_mem[16'h2237] <= 0;
        weight_mem[16'h2238] <= 0;
        weight_mem[16'h2239] <= 0;
        weight_mem[16'h223A] <= 0;
        weight_mem[16'h223B] <= 0;
        weight_mem[16'h223C] <= 0;
        weight_mem[16'h223D] <= 0;
        weight_mem[16'h223E] <= 0;
        weight_mem[16'h223F] <= 0;
        weight_mem[16'h2240] <= 0;
        weight_mem[16'h2241] <= 0;
        weight_mem[16'h2242] <= 0;
        weight_mem[16'h2243] <= 0;
        weight_mem[16'h2244] <= 0;
        weight_mem[16'h2245] <= 0;
        weight_mem[16'h2246] <= 0;
        weight_mem[16'h2247] <= 0;
        weight_mem[16'h2248] <= 0;
        weight_mem[16'h2249] <= 0;
        weight_mem[16'h224A] <= 0;
        weight_mem[16'h224B] <= 0;
        weight_mem[16'h224C] <= 0;
        weight_mem[16'h224D] <= 0;
        weight_mem[16'h224E] <= 0;
        weight_mem[16'h224F] <= 0;
        weight_mem[16'h2250] <= 0;
        weight_mem[16'h2251] <= 0;
        weight_mem[16'h2252] <= 0;
        weight_mem[16'h2253] <= 0;
        weight_mem[16'h2254] <= 0;
        weight_mem[16'h2255] <= 0;
        weight_mem[16'h2256] <= 0;
        weight_mem[16'h2257] <= 0;
        weight_mem[16'h2258] <= 0;
        weight_mem[16'h2259] <= 0;
        weight_mem[16'h225A] <= 0;
        weight_mem[16'h225B] <= 0;
        weight_mem[16'h225C] <= 0;
        weight_mem[16'h225D] <= 0;
        weight_mem[16'h225E] <= 0;
        weight_mem[16'h225F] <= 0;
        weight_mem[16'h2260] <= 0;
        weight_mem[16'h2261] <= 0;
        weight_mem[16'h2262] <= 0;
        weight_mem[16'h2263] <= 0;
        weight_mem[16'h2264] <= 0;
        weight_mem[16'h2265] <= 0;
        weight_mem[16'h2266] <= 0;
        weight_mem[16'h2267] <= 0;
        weight_mem[16'h2268] <= 0;
        weight_mem[16'h2269] <= 0;
        weight_mem[16'h226A] <= 0;
        weight_mem[16'h226B] <= 0;
        weight_mem[16'h226C] <= 0;
        weight_mem[16'h226D] <= 0;
        weight_mem[16'h226E] <= 0;
        weight_mem[16'h226F] <= 0;
        weight_mem[16'h2270] <= 0;
        weight_mem[16'h2271] <= 0;
        weight_mem[16'h2272] <= 0;
        weight_mem[16'h2273] <= 0;
        weight_mem[16'h2274] <= 0;
        weight_mem[16'h2275] <= 0;
        weight_mem[16'h2276] <= 0;
        weight_mem[16'h2277] <= 0;
        weight_mem[16'h2278] <= 0;
        weight_mem[16'h2279] <= 0;
        weight_mem[16'h227A] <= 0;
        weight_mem[16'h227B] <= 0;
        weight_mem[16'h227C] <= 0;
        weight_mem[16'h227D] <= 0;
        weight_mem[16'h227E] <= 0;
        weight_mem[16'h227F] <= 0;
        weight_mem[16'h2280] <= 0;
        weight_mem[16'h2281] <= 0;
        weight_mem[16'h2282] <= 0;
        weight_mem[16'h2283] <= 0;
        weight_mem[16'h2284] <= 0;
        weight_mem[16'h2285] <= 0;
        weight_mem[16'h2286] <= 0;
        weight_mem[16'h2287] <= 0;
        weight_mem[16'h2288] <= 0;
        weight_mem[16'h2289] <= 0;
        weight_mem[16'h228A] <= 0;
        weight_mem[16'h228B] <= 0;
        weight_mem[16'h228C] <= 0;
        weight_mem[16'h228D] <= 0;
        weight_mem[16'h228E] <= 0;
        weight_mem[16'h228F] <= 0;
        weight_mem[16'h2290] <= 0;
        weight_mem[16'h2291] <= 0;
        weight_mem[16'h2292] <= 0;
        weight_mem[16'h2293] <= 0;
        weight_mem[16'h2294] <= 0;
        weight_mem[16'h2295] <= 0;
        weight_mem[16'h2296] <= 0;
        weight_mem[16'h2297] <= 0;
        weight_mem[16'h2298] <= 0;
        weight_mem[16'h2299] <= 0;
        weight_mem[16'h229A] <= 0;
        weight_mem[16'h229B] <= 0;
        weight_mem[16'h229C] <= 0;
        weight_mem[16'h229D] <= 0;
        weight_mem[16'h229E] <= 0;
        weight_mem[16'h229F] <= 0;
        weight_mem[16'h22A0] <= 0;
        weight_mem[16'h22A1] <= 0;
        weight_mem[16'h22A2] <= 0;
        weight_mem[16'h22A3] <= 0;
        weight_mem[16'h22A4] <= 0;
        weight_mem[16'h22A5] <= 0;
        weight_mem[16'h22A6] <= 0;
        weight_mem[16'h22A7] <= 0;
        weight_mem[16'h22A8] <= 0;
        weight_mem[16'h22A9] <= 0;
        weight_mem[16'h22AA] <= 0;
        weight_mem[16'h22AB] <= 0;
        weight_mem[16'h22AC] <= 0;
        weight_mem[16'h22AD] <= 0;
        weight_mem[16'h22AE] <= 0;
        weight_mem[16'h22AF] <= 0;
        weight_mem[16'h22B0] <= 0;
        weight_mem[16'h22B1] <= 0;
        weight_mem[16'h22B2] <= 0;
        weight_mem[16'h22B3] <= 0;
        weight_mem[16'h22B4] <= 0;
        weight_mem[16'h22B5] <= 0;
        weight_mem[16'h22B6] <= 0;
        weight_mem[16'h22B7] <= 0;
        weight_mem[16'h22B8] <= 0;
        weight_mem[16'h22B9] <= 0;
        weight_mem[16'h22BA] <= 0;
        weight_mem[16'h22BB] <= 0;
        weight_mem[16'h22BC] <= 0;
        weight_mem[16'h22BD] <= 0;
        weight_mem[16'h22BE] <= 0;
        weight_mem[16'h22BF] <= 0;
        weight_mem[16'h22C0] <= 0;
        weight_mem[16'h22C1] <= 0;
        weight_mem[16'h22C2] <= 0;
        weight_mem[16'h22C3] <= 0;
        weight_mem[16'h22C4] <= 0;
        weight_mem[16'h22C5] <= 0;
        weight_mem[16'h22C6] <= 0;
        weight_mem[16'h22C7] <= 0;
        weight_mem[16'h22C8] <= 0;
        weight_mem[16'h22C9] <= 0;
        weight_mem[16'h22CA] <= 0;
        weight_mem[16'h22CB] <= 0;
        weight_mem[16'h22CC] <= 0;
        weight_mem[16'h22CD] <= 0;
        weight_mem[16'h22CE] <= 0;
        weight_mem[16'h22CF] <= 0;
        weight_mem[16'h22D0] <= 0;
        weight_mem[16'h22D1] <= 0;
        weight_mem[16'h22D2] <= 0;
        weight_mem[16'h22D3] <= 0;
        weight_mem[16'h22D4] <= 0;
        weight_mem[16'h22D5] <= 0;
        weight_mem[16'h22D6] <= 0;
        weight_mem[16'h22D7] <= 0;
        weight_mem[16'h22D8] <= 0;
        weight_mem[16'h22D9] <= 0;
        weight_mem[16'h22DA] <= 0;
        weight_mem[16'h22DB] <= 0;
        weight_mem[16'h22DC] <= 0;
        weight_mem[16'h22DD] <= 0;
        weight_mem[16'h22DE] <= 0;
        weight_mem[16'h22DF] <= 0;
        weight_mem[16'h22E0] <= 0;
        weight_mem[16'h22E1] <= 0;
        weight_mem[16'h22E2] <= 0;
        weight_mem[16'h22E3] <= 0;
        weight_mem[16'h22E4] <= 0;
        weight_mem[16'h22E5] <= 0;
        weight_mem[16'h22E6] <= 0;
        weight_mem[16'h22E7] <= 0;
        weight_mem[16'h22E8] <= 0;
        weight_mem[16'h22E9] <= 0;
        weight_mem[16'h22EA] <= 0;
        weight_mem[16'h22EB] <= 0;
        weight_mem[16'h22EC] <= 0;
        weight_mem[16'h22ED] <= 0;
        weight_mem[16'h22EE] <= 0;
        weight_mem[16'h22EF] <= 0;
        weight_mem[16'h22F0] <= 0;
        weight_mem[16'h22F1] <= 0;
        weight_mem[16'h22F2] <= 0;
        weight_mem[16'h22F3] <= 0;
        weight_mem[16'h22F4] <= 0;
        weight_mem[16'h22F5] <= 0;
        weight_mem[16'h22F6] <= 0;
        weight_mem[16'h22F7] <= 0;
        weight_mem[16'h22F8] <= 0;
        weight_mem[16'h22F9] <= 0;
        weight_mem[16'h22FA] <= 0;
        weight_mem[16'h22FB] <= 0;
        weight_mem[16'h22FC] <= 0;
        weight_mem[16'h22FD] <= 0;
        weight_mem[16'h22FE] <= 0;
        weight_mem[16'h22FF] <= 0;
        weight_mem[16'h2300] <= 0;
        weight_mem[16'h2301] <= 0;
        weight_mem[16'h2302] <= 0;
        weight_mem[16'h2303] <= 0;
        weight_mem[16'h2304] <= 0;
        weight_mem[16'h2305] <= 0;
        weight_mem[16'h2306] <= 0;
        weight_mem[16'h2307] <= 0;
        weight_mem[16'h2308] <= 0;
        weight_mem[16'h2309] <= 0;
        weight_mem[16'h230A] <= 0;
        weight_mem[16'h230B] <= 0;
        weight_mem[16'h230C] <= 0;
        weight_mem[16'h230D] <= 0;
        weight_mem[16'h230E] <= 0;
        weight_mem[16'h230F] <= 0;
        weight_mem[16'h2310] <= 0;
        weight_mem[16'h2311] <= 0;
        weight_mem[16'h2312] <= 0;
        weight_mem[16'h2313] <= 0;
        weight_mem[16'h2314] <= 0;
        weight_mem[16'h2315] <= 0;
        weight_mem[16'h2316] <= 0;
        weight_mem[16'h2317] <= 0;
        weight_mem[16'h2318] <= 0;
        weight_mem[16'h2319] <= 0;
        weight_mem[16'h231A] <= 0;
        weight_mem[16'h231B] <= 0;
        weight_mem[16'h231C] <= 0;
        weight_mem[16'h231D] <= 0;
        weight_mem[16'h231E] <= 0;
        weight_mem[16'h231F] <= 0;
        weight_mem[16'h2320] <= 0;
        weight_mem[16'h2321] <= 0;
        weight_mem[16'h2322] <= 0;
        weight_mem[16'h2323] <= 0;
        weight_mem[16'h2324] <= 0;
        weight_mem[16'h2325] <= 0;
        weight_mem[16'h2326] <= 0;
        weight_mem[16'h2327] <= 0;
        weight_mem[16'h2328] <= 0;
        weight_mem[16'h2329] <= 0;
        weight_mem[16'h232A] <= 0;
        weight_mem[16'h232B] <= 0;
        weight_mem[16'h232C] <= 0;
        weight_mem[16'h232D] <= 0;
        weight_mem[16'h232E] <= 0;
        weight_mem[16'h232F] <= 0;
        weight_mem[16'h2330] <= 0;
        weight_mem[16'h2331] <= 0;
        weight_mem[16'h2332] <= 0;
        weight_mem[16'h2333] <= 0;
        weight_mem[16'h2334] <= 0;
        weight_mem[16'h2335] <= 0;
        weight_mem[16'h2336] <= 0;
        weight_mem[16'h2337] <= 0;
        weight_mem[16'h2338] <= 0;
        weight_mem[16'h2339] <= 0;
        weight_mem[16'h233A] <= 0;
        weight_mem[16'h233B] <= 0;
        weight_mem[16'h233C] <= 0;
        weight_mem[16'h233D] <= 0;
        weight_mem[16'h233E] <= 0;
        weight_mem[16'h233F] <= 0;
        weight_mem[16'h2340] <= 0;
        weight_mem[16'h2341] <= 0;
        weight_mem[16'h2342] <= 0;
        weight_mem[16'h2343] <= 0;
        weight_mem[16'h2344] <= 0;
        weight_mem[16'h2345] <= 0;
        weight_mem[16'h2346] <= 0;
        weight_mem[16'h2347] <= 0;
        weight_mem[16'h2348] <= 0;
        weight_mem[16'h2349] <= 0;
        weight_mem[16'h234A] <= 0;
        weight_mem[16'h234B] <= 0;
        weight_mem[16'h234C] <= 0;
        weight_mem[16'h234D] <= 0;
        weight_mem[16'h234E] <= 0;
        weight_mem[16'h234F] <= 0;
        weight_mem[16'h2350] <= 0;
        weight_mem[16'h2351] <= 0;
        weight_mem[16'h2352] <= 0;
        weight_mem[16'h2353] <= 0;
        weight_mem[16'h2354] <= 0;
        weight_mem[16'h2355] <= 0;
        weight_mem[16'h2356] <= 0;
        weight_mem[16'h2357] <= 0;
        weight_mem[16'h2358] <= 0;
        weight_mem[16'h2359] <= 0;
        weight_mem[16'h235A] <= 0;
        weight_mem[16'h235B] <= 0;
        weight_mem[16'h235C] <= 0;
        weight_mem[16'h235D] <= 0;
        weight_mem[16'h235E] <= 0;
        weight_mem[16'h235F] <= 0;
        weight_mem[16'h2360] <= 0;
        weight_mem[16'h2361] <= 0;
        weight_mem[16'h2362] <= 0;
        weight_mem[16'h2363] <= 0;
        weight_mem[16'h2364] <= 0;
        weight_mem[16'h2365] <= 0;
        weight_mem[16'h2366] <= 0;
        weight_mem[16'h2367] <= 0;
        weight_mem[16'h2368] <= 0;
        weight_mem[16'h2369] <= 0;
        weight_mem[16'h236A] <= 0;
        weight_mem[16'h236B] <= 0;
        weight_mem[16'h236C] <= 0;
        weight_mem[16'h236D] <= 0;
        weight_mem[16'h236E] <= 0;
        weight_mem[16'h236F] <= 0;
        weight_mem[16'h2370] <= 0;
        weight_mem[16'h2371] <= 0;
        weight_mem[16'h2372] <= 0;
        weight_mem[16'h2373] <= 0;
        weight_mem[16'h2374] <= 0;
        weight_mem[16'h2375] <= 0;
        weight_mem[16'h2376] <= 0;
        weight_mem[16'h2377] <= 0;
        weight_mem[16'h2378] <= 0;
        weight_mem[16'h2379] <= 0;
        weight_mem[16'h237A] <= 0;
        weight_mem[16'h237B] <= 0;
        weight_mem[16'h237C] <= 0;
        weight_mem[16'h237D] <= 0;
        weight_mem[16'h237E] <= 0;
        weight_mem[16'h237F] <= 0;
        weight_mem[16'h2380] <= 0;
        weight_mem[16'h2381] <= 0;
        weight_mem[16'h2382] <= 0;
        weight_mem[16'h2383] <= 0;
        weight_mem[16'h2384] <= 0;
        weight_mem[16'h2385] <= 0;
        weight_mem[16'h2386] <= 0;
        weight_mem[16'h2387] <= 0;
        weight_mem[16'h2388] <= 0;
        weight_mem[16'h2389] <= 0;
        weight_mem[16'h238A] <= 0;
        weight_mem[16'h238B] <= 0;
        weight_mem[16'h238C] <= 0;
        weight_mem[16'h238D] <= 0;
        weight_mem[16'h238E] <= 0;
        weight_mem[16'h238F] <= 0;
        weight_mem[16'h2390] <= 0;
        weight_mem[16'h2391] <= 0;
        weight_mem[16'h2392] <= 0;
        weight_mem[16'h2393] <= 0;
        weight_mem[16'h2394] <= 0;
        weight_mem[16'h2395] <= 0;
        weight_mem[16'h2396] <= 0;
        weight_mem[16'h2397] <= 0;
        weight_mem[16'h2398] <= 0;
        weight_mem[16'h2399] <= 0;
        weight_mem[16'h239A] <= 0;
        weight_mem[16'h239B] <= 0;
        weight_mem[16'h239C] <= 0;
        weight_mem[16'h239D] <= 0;
        weight_mem[16'h239E] <= 0;
        weight_mem[16'h239F] <= 0;
        weight_mem[16'h23A0] <= 0;
        weight_mem[16'h23A1] <= 0;
        weight_mem[16'h23A2] <= 0;
        weight_mem[16'h23A3] <= 0;
        weight_mem[16'h23A4] <= 0;
        weight_mem[16'h23A5] <= 0;
        weight_mem[16'h23A6] <= 0;
        weight_mem[16'h23A7] <= 0;
        weight_mem[16'h23A8] <= 0;
        weight_mem[16'h23A9] <= 0;
        weight_mem[16'h23AA] <= 0;
        weight_mem[16'h23AB] <= 0;
        weight_mem[16'h23AC] <= 0;
        weight_mem[16'h23AD] <= 0;
        weight_mem[16'h23AE] <= 0;
        weight_mem[16'h23AF] <= 0;

        // layer 1 neuron 18
        weight_mem[16'h2400] <= 0;
        weight_mem[16'h2401] <= 0;
        weight_mem[16'h2402] <= 0;
        weight_mem[16'h2403] <= 0;
        weight_mem[16'h2404] <= 0;
        weight_mem[16'h2405] <= 0;
        weight_mem[16'h2406] <= 0;
        weight_mem[16'h2407] <= 0;
        weight_mem[16'h2408] <= 0;
        weight_mem[16'h2409] <= 0;
        weight_mem[16'h240A] <= 0;
        weight_mem[16'h240B] <= 0;
        weight_mem[16'h240C] <= 0;
        weight_mem[16'h240D] <= 0;
        weight_mem[16'h240E] <= 0;
        weight_mem[16'h240F] <= 0;
        weight_mem[16'h2410] <= 0;
        weight_mem[16'h2411] <= 0;
        weight_mem[16'h2412] <= 0;
        weight_mem[16'h2413] <= 0;
        weight_mem[16'h2414] <= 0;
        weight_mem[16'h2415] <= 0;
        weight_mem[16'h2416] <= 0;
        weight_mem[16'h2417] <= 0;
        weight_mem[16'h2418] <= 0;
        weight_mem[16'h2419] <= 0;
        weight_mem[16'h241A] <= 0;
        weight_mem[16'h241B] <= 0;
        weight_mem[16'h241C] <= 0;
        weight_mem[16'h241D] <= 0;
        weight_mem[16'h241E] <= 0;
        weight_mem[16'h241F] <= 0;
        weight_mem[16'h2420] <= 0;
        weight_mem[16'h2421] <= 0;
        weight_mem[16'h2422] <= 0;
        weight_mem[16'h2423] <= 0;
        weight_mem[16'h2424] <= 0;
        weight_mem[16'h2425] <= 0;
        weight_mem[16'h2426] <= 0;
        weight_mem[16'h2427] <= 0;
        weight_mem[16'h2428] <= 0;
        weight_mem[16'h2429] <= 0;
        weight_mem[16'h242A] <= 0;
        weight_mem[16'h242B] <= 0;
        weight_mem[16'h242C] <= 0;
        weight_mem[16'h242D] <= 0;
        weight_mem[16'h242E] <= 0;
        weight_mem[16'h242F] <= 0;
        weight_mem[16'h2430] <= 0;
        weight_mem[16'h2431] <= 0;
        weight_mem[16'h2432] <= 0;
        weight_mem[16'h2433] <= 0;
        weight_mem[16'h2434] <= 0;
        weight_mem[16'h2435] <= 0;
        weight_mem[16'h2436] <= 0;
        weight_mem[16'h2437] <= 0;
        weight_mem[16'h2438] <= 0;
        weight_mem[16'h2439] <= 0;
        weight_mem[16'h243A] <= 0;
        weight_mem[16'h243B] <= 0;
        weight_mem[16'h243C] <= 0;
        weight_mem[16'h243D] <= 0;
        weight_mem[16'h243E] <= 0;
        weight_mem[16'h243F] <= 0;
        weight_mem[16'h2440] <= 0;
        weight_mem[16'h2441] <= 0;
        weight_mem[16'h2442] <= 0;
        weight_mem[16'h2443] <= 0;
        weight_mem[16'h2444] <= 0;
        weight_mem[16'h2445] <= 0;
        weight_mem[16'h2446] <= 0;
        weight_mem[16'h2447] <= 0;
        weight_mem[16'h2448] <= 0;
        weight_mem[16'h2449] <= 0;
        weight_mem[16'h244A] <= 0;
        weight_mem[16'h244B] <= 0;
        weight_mem[16'h244C] <= 0;
        weight_mem[16'h244D] <= 0;
        weight_mem[16'h244E] <= 0;
        weight_mem[16'h244F] <= 0;
        weight_mem[16'h2450] <= 0;
        weight_mem[16'h2451] <= 0;
        weight_mem[16'h2452] <= 0;
        weight_mem[16'h2453] <= 0;
        weight_mem[16'h2454] <= 0;
        weight_mem[16'h2455] <= 0;
        weight_mem[16'h2456] <= 0;
        weight_mem[16'h2457] <= 0;
        weight_mem[16'h2458] <= 0;
        weight_mem[16'h2459] <= 0;
        weight_mem[16'h245A] <= 0;
        weight_mem[16'h245B] <= 0;
        weight_mem[16'h245C] <= 0;
        weight_mem[16'h245D] <= 0;
        weight_mem[16'h245E] <= 0;
        weight_mem[16'h245F] <= 0;
        weight_mem[16'h2460] <= 0;
        weight_mem[16'h2461] <= 0;
        weight_mem[16'h2462] <= 0;
        weight_mem[16'h2463] <= 0;
        weight_mem[16'h2464] <= 0;
        weight_mem[16'h2465] <= 0;
        weight_mem[16'h2466] <= 0;
        weight_mem[16'h2467] <= 0;
        weight_mem[16'h2468] <= 0;
        weight_mem[16'h2469] <= 0;
        weight_mem[16'h246A] <= 0;
        weight_mem[16'h246B] <= 0;
        weight_mem[16'h246C] <= 0;
        weight_mem[16'h246D] <= 0;
        weight_mem[16'h246E] <= 0;
        weight_mem[16'h246F] <= 0;
        weight_mem[16'h2470] <= 0;
        weight_mem[16'h2471] <= 0;
        weight_mem[16'h2472] <= 0;
        weight_mem[16'h2473] <= 0;
        weight_mem[16'h2474] <= 0;
        weight_mem[16'h2475] <= 0;
        weight_mem[16'h2476] <= 0;
        weight_mem[16'h2477] <= 0;
        weight_mem[16'h2478] <= 0;
        weight_mem[16'h2479] <= 0;
        weight_mem[16'h247A] <= 0;
        weight_mem[16'h247B] <= 0;
        weight_mem[16'h247C] <= 0;
        weight_mem[16'h247D] <= 0;
        weight_mem[16'h247E] <= 0;
        weight_mem[16'h247F] <= 0;
        weight_mem[16'h2480] <= 0;
        weight_mem[16'h2481] <= 0;
        weight_mem[16'h2482] <= 0;
        weight_mem[16'h2483] <= 0;
        weight_mem[16'h2484] <= 0;
        weight_mem[16'h2485] <= 0;
        weight_mem[16'h2486] <= 0;
        weight_mem[16'h2487] <= 0;
        weight_mem[16'h2488] <= 0;
        weight_mem[16'h2489] <= 0;
        weight_mem[16'h248A] <= 0;
        weight_mem[16'h248B] <= 0;
        weight_mem[16'h248C] <= 0;
        weight_mem[16'h248D] <= 0;
        weight_mem[16'h248E] <= 0;
        weight_mem[16'h248F] <= 0;
        weight_mem[16'h2490] <= 0;
        weight_mem[16'h2491] <= 0;
        weight_mem[16'h2492] <= 0;
        weight_mem[16'h2493] <= 0;
        weight_mem[16'h2494] <= 0;
        weight_mem[16'h2495] <= 0;
        weight_mem[16'h2496] <= 0;
        weight_mem[16'h2497] <= 0;
        weight_mem[16'h2498] <= 0;
        weight_mem[16'h2499] <= 0;
        weight_mem[16'h249A] <= 0;
        weight_mem[16'h249B] <= 0;
        weight_mem[16'h249C] <= 0;
        weight_mem[16'h249D] <= 0;
        weight_mem[16'h249E] <= 0;
        weight_mem[16'h249F] <= 0;
        weight_mem[16'h24A0] <= 0;
        weight_mem[16'h24A1] <= 0;
        weight_mem[16'h24A2] <= 0;
        weight_mem[16'h24A3] <= 0;
        weight_mem[16'h24A4] <= 0;
        weight_mem[16'h24A5] <= 0;
        weight_mem[16'h24A6] <= 0;
        weight_mem[16'h24A7] <= 0;
        weight_mem[16'h24A8] <= 0;
        weight_mem[16'h24A9] <= 0;
        weight_mem[16'h24AA] <= 0;
        weight_mem[16'h24AB] <= 0;
        weight_mem[16'h24AC] <= 0;
        weight_mem[16'h24AD] <= 0;
        weight_mem[16'h24AE] <= 0;
        weight_mem[16'h24AF] <= 0;
        weight_mem[16'h24B0] <= 0;
        weight_mem[16'h24B1] <= 0;
        weight_mem[16'h24B2] <= 0;
        weight_mem[16'h24B3] <= 0;
        weight_mem[16'h24B4] <= 0;
        weight_mem[16'h24B5] <= 0;
        weight_mem[16'h24B6] <= 0;
        weight_mem[16'h24B7] <= 0;
        weight_mem[16'h24B8] <= 0;
        weight_mem[16'h24B9] <= 0;
        weight_mem[16'h24BA] <= 0;
        weight_mem[16'h24BB] <= 0;
        weight_mem[16'h24BC] <= 0;
        weight_mem[16'h24BD] <= 0;
        weight_mem[16'h24BE] <= 0;
        weight_mem[16'h24BF] <= 0;
        weight_mem[16'h24C0] <= 0;
        weight_mem[16'h24C1] <= 0;
        weight_mem[16'h24C2] <= 0;
        weight_mem[16'h24C3] <= 0;
        weight_mem[16'h24C4] <= 0;
        weight_mem[16'h24C5] <= 0;
        weight_mem[16'h24C6] <= 0;
        weight_mem[16'h24C7] <= 0;
        weight_mem[16'h24C8] <= 0;
        weight_mem[16'h24C9] <= 0;
        weight_mem[16'h24CA] <= 0;
        weight_mem[16'h24CB] <= 0;
        weight_mem[16'h24CC] <= 0;
        weight_mem[16'h24CD] <= 0;
        weight_mem[16'h24CE] <= 0;
        weight_mem[16'h24CF] <= 0;
        weight_mem[16'h24D0] <= 0;
        weight_mem[16'h24D1] <= 0;
        weight_mem[16'h24D2] <= 0;
        weight_mem[16'h24D3] <= 0;
        weight_mem[16'h24D4] <= 0;
        weight_mem[16'h24D5] <= 0;
        weight_mem[16'h24D6] <= 0;
        weight_mem[16'h24D7] <= 0;
        weight_mem[16'h24D8] <= 0;
        weight_mem[16'h24D9] <= 0;
        weight_mem[16'h24DA] <= 0;
        weight_mem[16'h24DB] <= 0;
        weight_mem[16'h24DC] <= 0;
        weight_mem[16'h24DD] <= 0;
        weight_mem[16'h24DE] <= 0;
        weight_mem[16'h24DF] <= 0;
        weight_mem[16'h24E0] <= 0;
        weight_mem[16'h24E1] <= 0;
        weight_mem[16'h24E2] <= 0;
        weight_mem[16'h24E3] <= 0;
        weight_mem[16'h24E4] <= 0;
        weight_mem[16'h24E5] <= 0;
        weight_mem[16'h24E6] <= 0;
        weight_mem[16'h24E7] <= 0;
        weight_mem[16'h24E8] <= 0;
        weight_mem[16'h24E9] <= 0;
        weight_mem[16'h24EA] <= 0;
        weight_mem[16'h24EB] <= 0;
        weight_mem[16'h24EC] <= 0;
        weight_mem[16'h24ED] <= 0;
        weight_mem[16'h24EE] <= 0;
        weight_mem[16'h24EF] <= 0;
        weight_mem[16'h24F0] <= 0;
        weight_mem[16'h24F1] <= 0;
        weight_mem[16'h24F2] <= 0;
        weight_mem[16'h24F3] <= 0;
        weight_mem[16'h24F4] <= 0;
        weight_mem[16'h24F5] <= 0;
        weight_mem[16'h24F6] <= 0;
        weight_mem[16'h24F7] <= 0;
        weight_mem[16'h24F8] <= 0;
        weight_mem[16'h24F9] <= 0;
        weight_mem[16'h24FA] <= 0;
        weight_mem[16'h24FB] <= 0;
        weight_mem[16'h24FC] <= 0;
        weight_mem[16'h24FD] <= 0;
        weight_mem[16'h24FE] <= 0;
        weight_mem[16'h24FF] <= 0;
        weight_mem[16'h2500] <= 0;
        weight_mem[16'h2501] <= 0;
        weight_mem[16'h2502] <= 0;
        weight_mem[16'h2503] <= 0;
        weight_mem[16'h2504] <= 0;
        weight_mem[16'h2505] <= 0;
        weight_mem[16'h2506] <= 0;
        weight_mem[16'h2507] <= 0;
        weight_mem[16'h2508] <= 0;
        weight_mem[16'h2509] <= 0;
        weight_mem[16'h250A] <= 0;
        weight_mem[16'h250B] <= 0;
        weight_mem[16'h250C] <= 0;
        weight_mem[16'h250D] <= 0;
        weight_mem[16'h250E] <= 0;
        weight_mem[16'h250F] <= 0;
        weight_mem[16'h2510] <= 0;
        weight_mem[16'h2511] <= 0;
        weight_mem[16'h2512] <= 0;
        weight_mem[16'h2513] <= 0;
        weight_mem[16'h2514] <= 0;
        weight_mem[16'h2515] <= 0;
        weight_mem[16'h2516] <= 0;
        weight_mem[16'h2517] <= 0;
        weight_mem[16'h2518] <= 0;
        weight_mem[16'h2519] <= 0;
        weight_mem[16'h251A] <= 0;
        weight_mem[16'h251B] <= 0;
        weight_mem[16'h251C] <= 0;
        weight_mem[16'h251D] <= 0;
        weight_mem[16'h251E] <= 0;
        weight_mem[16'h251F] <= 0;
        weight_mem[16'h2520] <= 0;
        weight_mem[16'h2521] <= 0;
        weight_mem[16'h2522] <= 0;
        weight_mem[16'h2523] <= 0;
        weight_mem[16'h2524] <= 0;
        weight_mem[16'h2525] <= 0;
        weight_mem[16'h2526] <= 0;
        weight_mem[16'h2527] <= 0;
        weight_mem[16'h2528] <= 0;
        weight_mem[16'h2529] <= 0;
        weight_mem[16'h252A] <= 0;
        weight_mem[16'h252B] <= 0;
        weight_mem[16'h252C] <= 0;
        weight_mem[16'h252D] <= 0;
        weight_mem[16'h252E] <= 0;
        weight_mem[16'h252F] <= 0;
        weight_mem[16'h2530] <= 0;
        weight_mem[16'h2531] <= 0;
        weight_mem[16'h2532] <= 0;
        weight_mem[16'h2533] <= 0;
        weight_mem[16'h2534] <= 0;
        weight_mem[16'h2535] <= 0;
        weight_mem[16'h2536] <= 0;
        weight_mem[16'h2537] <= 0;
        weight_mem[16'h2538] <= 0;
        weight_mem[16'h2539] <= 0;
        weight_mem[16'h253A] <= 0;
        weight_mem[16'h253B] <= 0;
        weight_mem[16'h253C] <= 0;
        weight_mem[16'h253D] <= 0;
        weight_mem[16'h253E] <= 0;
        weight_mem[16'h253F] <= 0;
        weight_mem[16'h2540] <= 0;
        weight_mem[16'h2541] <= 0;
        weight_mem[16'h2542] <= 0;
        weight_mem[16'h2543] <= 0;
        weight_mem[16'h2544] <= 0;
        weight_mem[16'h2545] <= 0;
        weight_mem[16'h2546] <= 0;
        weight_mem[16'h2547] <= 0;
        weight_mem[16'h2548] <= 0;
        weight_mem[16'h2549] <= 0;
        weight_mem[16'h254A] <= 0;
        weight_mem[16'h254B] <= 0;
        weight_mem[16'h254C] <= 0;
        weight_mem[16'h254D] <= 0;
        weight_mem[16'h254E] <= 0;
        weight_mem[16'h254F] <= 0;
        weight_mem[16'h2550] <= 0;
        weight_mem[16'h2551] <= 0;
        weight_mem[16'h2552] <= 0;
        weight_mem[16'h2553] <= 0;
        weight_mem[16'h2554] <= 0;
        weight_mem[16'h2555] <= 0;
        weight_mem[16'h2556] <= 0;
        weight_mem[16'h2557] <= 0;
        weight_mem[16'h2558] <= 0;
        weight_mem[16'h2559] <= 0;
        weight_mem[16'h255A] <= 0;
        weight_mem[16'h255B] <= 0;
        weight_mem[16'h255C] <= 0;
        weight_mem[16'h255D] <= 0;
        weight_mem[16'h255E] <= 0;
        weight_mem[16'h255F] <= 0;
        weight_mem[16'h2560] <= 0;
        weight_mem[16'h2561] <= 0;
        weight_mem[16'h2562] <= 0;
        weight_mem[16'h2563] <= 0;
        weight_mem[16'h2564] <= 0;
        weight_mem[16'h2565] <= 0;
        weight_mem[16'h2566] <= 0;
        weight_mem[16'h2567] <= 0;
        weight_mem[16'h2568] <= 0;
        weight_mem[16'h2569] <= 0;
        weight_mem[16'h256A] <= 0;
        weight_mem[16'h256B] <= 0;
        weight_mem[16'h256C] <= 0;
        weight_mem[16'h256D] <= 0;
        weight_mem[16'h256E] <= 0;
        weight_mem[16'h256F] <= 0;
        weight_mem[16'h2570] <= 0;
        weight_mem[16'h2571] <= 0;
        weight_mem[16'h2572] <= 0;
        weight_mem[16'h2573] <= 0;
        weight_mem[16'h2574] <= 0;
        weight_mem[16'h2575] <= 0;
        weight_mem[16'h2576] <= 0;
        weight_mem[16'h2577] <= 0;
        weight_mem[16'h2578] <= 0;
        weight_mem[16'h2579] <= 0;
        weight_mem[16'h257A] <= 0;
        weight_mem[16'h257B] <= 0;
        weight_mem[16'h257C] <= 0;
        weight_mem[16'h257D] <= 0;
        weight_mem[16'h257E] <= 0;
        weight_mem[16'h257F] <= 0;
        weight_mem[16'h2580] <= 0;
        weight_mem[16'h2581] <= 0;
        weight_mem[16'h2582] <= 0;
        weight_mem[16'h2583] <= 0;
        weight_mem[16'h2584] <= 0;
        weight_mem[16'h2585] <= 0;
        weight_mem[16'h2586] <= 0;
        weight_mem[16'h2587] <= 0;
        weight_mem[16'h2588] <= 0;
        weight_mem[16'h2589] <= 0;
        weight_mem[16'h258A] <= 0;
        weight_mem[16'h258B] <= 0;
        weight_mem[16'h258C] <= 0;
        weight_mem[16'h258D] <= 0;
        weight_mem[16'h258E] <= 0;
        weight_mem[16'h258F] <= 0;
        weight_mem[16'h2590] <= 0;
        weight_mem[16'h2591] <= 0;
        weight_mem[16'h2592] <= 0;
        weight_mem[16'h2593] <= 0;
        weight_mem[16'h2594] <= 0;
        weight_mem[16'h2595] <= 0;
        weight_mem[16'h2596] <= 0;
        weight_mem[16'h2597] <= 0;
        weight_mem[16'h2598] <= 0;
        weight_mem[16'h2599] <= 0;
        weight_mem[16'h259A] <= 0;
        weight_mem[16'h259B] <= 0;
        weight_mem[16'h259C] <= 0;
        weight_mem[16'h259D] <= 0;
        weight_mem[16'h259E] <= 0;
        weight_mem[16'h259F] <= 0;
        weight_mem[16'h25A0] <= 0;
        weight_mem[16'h25A1] <= 0;
        weight_mem[16'h25A2] <= 0;
        weight_mem[16'h25A3] <= 0;
        weight_mem[16'h25A4] <= 0;
        weight_mem[16'h25A5] <= 0;
        weight_mem[16'h25A6] <= 0;
        weight_mem[16'h25A7] <= 0;
        weight_mem[16'h25A8] <= 0;
        weight_mem[16'h25A9] <= 0;
        weight_mem[16'h25AA] <= 0;
        weight_mem[16'h25AB] <= 0;
        weight_mem[16'h25AC] <= 0;
        weight_mem[16'h25AD] <= 0;
        weight_mem[16'h25AE] <= 0;
        weight_mem[16'h25AF] <= 0;

        // layer 1 neuron 19
        weight_mem[16'h2600] <= 0;
        weight_mem[16'h2601] <= 0;
        weight_mem[16'h2602] <= 0;
        weight_mem[16'h2603] <= 0;
        weight_mem[16'h2604] <= 0;
        weight_mem[16'h2605] <= 0;
        weight_mem[16'h2606] <= 0;
        weight_mem[16'h2607] <= 0;
        weight_mem[16'h2608] <= 0;
        weight_mem[16'h2609] <= 0;
        weight_mem[16'h260A] <= 0;
        weight_mem[16'h260B] <= 0;
        weight_mem[16'h260C] <= 0;
        weight_mem[16'h260D] <= 0;
        weight_mem[16'h260E] <= 0;
        weight_mem[16'h260F] <= 0;
        weight_mem[16'h2610] <= 0;
        weight_mem[16'h2611] <= 0;
        weight_mem[16'h2612] <= 0;
        weight_mem[16'h2613] <= 0;
        weight_mem[16'h2614] <= 0;
        weight_mem[16'h2615] <= 0;
        weight_mem[16'h2616] <= 0;
        weight_mem[16'h2617] <= 0;
        weight_mem[16'h2618] <= 0;
        weight_mem[16'h2619] <= 0;
        weight_mem[16'h261A] <= 0;
        weight_mem[16'h261B] <= 0;
        weight_mem[16'h261C] <= 0;
        weight_mem[16'h261D] <= 0;
        weight_mem[16'h261E] <= 0;
        weight_mem[16'h261F] <= 0;
        weight_mem[16'h2620] <= 0;
        weight_mem[16'h2621] <= 0;
        weight_mem[16'h2622] <= 0;
        weight_mem[16'h2623] <= 0;
        weight_mem[16'h2624] <= 0;
        weight_mem[16'h2625] <= 0;
        weight_mem[16'h2626] <= 0;
        weight_mem[16'h2627] <= 0;
        weight_mem[16'h2628] <= 0;
        weight_mem[16'h2629] <= 0;
        weight_mem[16'h262A] <= 0;
        weight_mem[16'h262B] <= 0;
        weight_mem[16'h262C] <= 0;
        weight_mem[16'h262D] <= 0;
        weight_mem[16'h262E] <= 0;
        weight_mem[16'h262F] <= 0;
        weight_mem[16'h2630] <= 0;
        weight_mem[16'h2631] <= 0;
        weight_mem[16'h2632] <= 0;
        weight_mem[16'h2633] <= 0;
        weight_mem[16'h2634] <= 0;
        weight_mem[16'h2635] <= 0;
        weight_mem[16'h2636] <= 0;
        weight_mem[16'h2637] <= 0;
        weight_mem[16'h2638] <= 0;
        weight_mem[16'h2639] <= 0;
        weight_mem[16'h263A] <= 0;
        weight_mem[16'h263B] <= 0;
        weight_mem[16'h263C] <= 0;
        weight_mem[16'h263D] <= 0;
        weight_mem[16'h263E] <= 0;
        weight_mem[16'h263F] <= 0;
        weight_mem[16'h2640] <= 0;
        weight_mem[16'h2641] <= 0;
        weight_mem[16'h2642] <= 0;
        weight_mem[16'h2643] <= 0;
        weight_mem[16'h2644] <= 0;
        weight_mem[16'h2645] <= 0;
        weight_mem[16'h2646] <= 0;
        weight_mem[16'h2647] <= 0;
        weight_mem[16'h2648] <= 0;
        weight_mem[16'h2649] <= 0;
        weight_mem[16'h264A] <= 0;
        weight_mem[16'h264B] <= 0;
        weight_mem[16'h264C] <= 0;
        weight_mem[16'h264D] <= 0;
        weight_mem[16'h264E] <= 0;
        weight_mem[16'h264F] <= 0;
        weight_mem[16'h2650] <= 0;
        weight_mem[16'h2651] <= 0;
        weight_mem[16'h2652] <= 0;
        weight_mem[16'h2653] <= 0;
        weight_mem[16'h2654] <= 0;
        weight_mem[16'h2655] <= 0;
        weight_mem[16'h2656] <= 0;
        weight_mem[16'h2657] <= 0;
        weight_mem[16'h2658] <= 0;
        weight_mem[16'h2659] <= 0;
        weight_mem[16'h265A] <= 0;
        weight_mem[16'h265B] <= 0;
        weight_mem[16'h265C] <= 0;
        weight_mem[16'h265D] <= 0;
        weight_mem[16'h265E] <= 0;
        weight_mem[16'h265F] <= 0;
        weight_mem[16'h2660] <= 0;
        weight_mem[16'h2661] <= 0;
        weight_mem[16'h2662] <= 0;
        weight_mem[16'h2663] <= 0;
        weight_mem[16'h2664] <= 0;
        weight_mem[16'h2665] <= 0;
        weight_mem[16'h2666] <= 0;
        weight_mem[16'h2667] <= 0;
        weight_mem[16'h2668] <= 0;
        weight_mem[16'h2669] <= 0;
        weight_mem[16'h266A] <= 0;
        weight_mem[16'h266B] <= 0;
        weight_mem[16'h266C] <= 0;
        weight_mem[16'h266D] <= 0;
        weight_mem[16'h266E] <= 0;
        weight_mem[16'h266F] <= 0;
        weight_mem[16'h2670] <= 0;
        weight_mem[16'h2671] <= 0;
        weight_mem[16'h2672] <= 0;
        weight_mem[16'h2673] <= 0;
        weight_mem[16'h2674] <= 0;
        weight_mem[16'h2675] <= 0;
        weight_mem[16'h2676] <= 0;
        weight_mem[16'h2677] <= 0;
        weight_mem[16'h2678] <= 0;
        weight_mem[16'h2679] <= 0;
        weight_mem[16'h267A] <= 0;
        weight_mem[16'h267B] <= 0;
        weight_mem[16'h267C] <= 0;
        weight_mem[16'h267D] <= 0;
        weight_mem[16'h267E] <= 0;
        weight_mem[16'h267F] <= 0;
        weight_mem[16'h2680] <= 0;
        weight_mem[16'h2681] <= 0;
        weight_mem[16'h2682] <= 0;
        weight_mem[16'h2683] <= 0;
        weight_mem[16'h2684] <= 0;
        weight_mem[16'h2685] <= 0;
        weight_mem[16'h2686] <= 0;
        weight_mem[16'h2687] <= 0;
        weight_mem[16'h2688] <= 0;
        weight_mem[16'h2689] <= 0;
        weight_mem[16'h268A] <= 0;
        weight_mem[16'h268B] <= 0;
        weight_mem[16'h268C] <= 0;
        weight_mem[16'h268D] <= 0;
        weight_mem[16'h268E] <= 0;
        weight_mem[16'h268F] <= 0;
        weight_mem[16'h2690] <= 0;
        weight_mem[16'h2691] <= 0;
        weight_mem[16'h2692] <= 0;
        weight_mem[16'h2693] <= 0;
        weight_mem[16'h2694] <= 0;
        weight_mem[16'h2695] <= 0;
        weight_mem[16'h2696] <= 0;
        weight_mem[16'h2697] <= 0;
        weight_mem[16'h2698] <= 0;
        weight_mem[16'h2699] <= 0;
        weight_mem[16'h269A] <= 0;
        weight_mem[16'h269B] <= 0;
        weight_mem[16'h269C] <= 0;
        weight_mem[16'h269D] <= 0;
        weight_mem[16'h269E] <= 0;
        weight_mem[16'h269F] <= 0;
        weight_mem[16'h26A0] <= 0;
        weight_mem[16'h26A1] <= 0;
        weight_mem[16'h26A2] <= 0;
        weight_mem[16'h26A3] <= 0;
        weight_mem[16'h26A4] <= 0;
        weight_mem[16'h26A5] <= 0;
        weight_mem[16'h26A6] <= 0;
        weight_mem[16'h26A7] <= 0;
        weight_mem[16'h26A8] <= 0;
        weight_mem[16'h26A9] <= 0;
        weight_mem[16'h26AA] <= 0;
        weight_mem[16'h26AB] <= 0;
        weight_mem[16'h26AC] <= 0;
        weight_mem[16'h26AD] <= 0;
        weight_mem[16'h26AE] <= 0;
        weight_mem[16'h26AF] <= 0;
        weight_mem[16'h26B0] <= 0;
        weight_mem[16'h26B1] <= 0;
        weight_mem[16'h26B2] <= 0;
        weight_mem[16'h26B3] <= 0;
        weight_mem[16'h26B4] <= 0;
        weight_mem[16'h26B5] <= 0;
        weight_mem[16'h26B6] <= 0;
        weight_mem[16'h26B7] <= 0;
        weight_mem[16'h26B8] <= 0;
        weight_mem[16'h26B9] <= 0;
        weight_mem[16'h26BA] <= 0;
        weight_mem[16'h26BB] <= 0;
        weight_mem[16'h26BC] <= 0;
        weight_mem[16'h26BD] <= 0;
        weight_mem[16'h26BE] <= 0;
        weight_mem[16'h26BF] <= 0;
        weight_mem[16'h26C0] <= 0;
        weight_mem[16'h26C1] <= 0;
        weight_mem[16'h26C2] <= 0;
        weight_mem[16'h26C3] <= 0;
        weight_mem[16'h26C4] <= 0;
        weight_mem[16'h26C5] <= 0;
        weight_mem[16'h26C6] <= 0;
        weight_mem[16'h26C7] <= 0;
        weight_mem[16'h26C8] <= 0;
        weight_mem[16'h26C9] <= 0;
        weight_mem[16'h26CA] <= 0;
        weight_mem[16'h26CB] <= 0;
        weight_mem[16'h26CC] <= 0;
        weight_mem[16'h26CD] <= 0;
        weight_mem[16'h26CE] <= 0;
        weight_mem[16'h26CF] <= 0;
        weight_mem[16'h26D0] <= 0;
        weight_mem[16'h26D1] <= 0;
        weight_mem[16'h26D2] <= 0;
        weight_mem[16'h26D3] <= 0;
        weight_mem[16'h26D4] <= 0;
        weight_mem[16'h26D5] <= 0;
        weight_mem[16'h26D6] <= 0;
        weight_mem[16'h26D7] <= 0;
        weight_mem[16'h26D8] <= 0;
        weight_mem[16'h26D9] <= 0;
        weight_mem[16'h26DA] <= 0;
        weight_mem[16'h26DB] <= 0;
        weight_mem[16'h26DC] <= 0;
        weight_mem[16'h26DD] <= 0;
        weight_mem[16'h26DE] <= 0;
        weight_mem[16'h26DF] <= 0;
        weight_mem[16'h26E0] <= 0;
        weight_mem[16'h26E1] <= 0;
        weight_mem[16'h26E2] <= 0;
        weight_mem[16'h26E3] <= 0;
        weight_mem[16'h26E4] <= 0;
        weight_mem[16'h26E5] <= 0;
        weight_mem[16'h26E6] <= 0;
        weight_mem[16'h26E7] <= 0;
        weight_mem[16'h26E8] <= 0;
        weight_mem[16'h26E9] <= 0;
        weight_mem[16'h26EA] <= 0;
        weight_mem[16'h26EB] <= 0;
        weight_mem[16'h26EC] <= 0;
        weight_mem[16'h26ED] <= 0;
        weight_mem[16'h26EE] <= 0;
        weight_mem[16'h26EF] <= 0;
        weight_mem[16'h26F0] <= 0;
        weight_mem[16'h26F1] <= 0;
        weight_mem[16'h26F2] <= 0;
        weight_mem[16'h26F3] <= 0;
        weight_mem[16'h26F4] <= 0;
        weight_mem[16'h26F5] <= 0;
        weight_mem[16'h26F6] <= 0;
        weight_mem[16'h26F7] <= 0;
        weight_mem[16'h26F8] <= 0;
        weight_mem[16'h26F9] <= 0;
        weight_mem[16'h26FA] <= 0;
        weight_mem[16'h26FB] <= 0;
        weight_mem[16'h26FC] <= 0;
        weight_mem[16'h26FD] <= 0;
        weight_mem[16'h26FE] <= 0;
        weight_mem[16'h26FF] <= 0;
        weight_mem[16'h2700] <= 0;
        weight_mem[16'h2701] <= 0;
        weight_mem[16'h2702] <= 0;
        weight_mem[16'h2703] <= 0;
        weight_mem[16'h2704] <= 0;
        weight_mem[16'h2705] <= 0;
        weight_mem[16'h2706] <= 0;
        weight_mem[16'h2707] <= 0;
        weight_mem[16'h2708] <= 0;
        weight_mem[16'h2709] <= 0;
        weight_mem[16'h270A] <= 0;
        weight_mem[16'h270B] <= 0;
        weight_mem[16'h270C] <= 0;
        weight_mem[16'h270D] <= 0;
        weight_mem[16'h270E] <= 0;
        weight_mem[16'h270F] <= 0;
        weight_mem[16'h2710] <= 0;
        weight_mem[16'h2711] <= 0;
        weight_mem[16'h2712] <= 0;
        weight_mem[16'h2713] <= 0;
        weight_mem[16'h2714] <= 0;
        weight_mem[16'h2715] <= 0;
        weight_mem[16'h2716] <= 0;
        weight_mem[16'h2717] <= 0;
        weight_mem[16'h2718] <= 0;
        weight_mem[16'h2719] <= 0;
        weight_mem[16'h271A] <= 0;
        weight_mem[16'h271B] <= 0;
        weight_mem[16'h271C] <= 0;
        weight_mem[16'h271D] <= 0;
        weight_mem[16'h271E] <= 0;
        weight_mem[16'h271F] <= 0;
        weight_mem[16'h2720] <= 0;
        weight_mem[16'h2721] <= 0;
        weight_mem[16'h2722] <= 0;
        weight_mem[16'h2723] <= 0;
        weight_mem[16'h2724] <= 0;
        weight_mem[16'h2725] <= 0;
        weight_mem[16'h2726] <= 0;
        weight_mem[16'h2727] <= 0;
        weight_mem[16'h2728] <= 0;
        weight_mem[16'h2729] <= 0;
        weight_mem[16'h272A] <= 0;
        weight_mem[16'h272B] <= 0;
        weight_mem[16'h272C] <= 0;
        weight_mem[16'h272D] <= 0;
        weight_mem[16'h272E] <= 0;
        weight_mem[16'h272F] <= 0;
        weight_mem[16'h2730] <= 0;
        weight_mem[16'h2731] <= 0;
        weight_mem[16'h2732] <= 0;
        weight_mem[16'h2733] <= 0;
        weight_mem[16'h2734] <= 0;
        weight_mem[16'h2735] <= 0;
        weight_mem[16'h2736] <= 0;
        weight_mem[16'h2737] <= 0;
        weight_mem[16'h2738] <= 0;
        weight_mem[16'h2739] <= 0;
        weight_mem[16'h273A] <= 0;
        weight_mem[16'h273B] <= 0;
        weight_mem[16'h273C] <= 0;
        weight_mem[16'h273D] <= 0;
        weight_mem[16'h273E] <= 0;
        weight_mem[16'h273F] <= 0;
        weight_mem[16'h2740] <= 0;
        weight_mem[16'h2741] <= 0;
        weight_mem[16'h2742] <= 0;
        weight_mem[16'h2743] <= 0;
        weight_mem[16'h2744] <= 0;
        weight_mem[16'h2745] <= 0;
        weight_mem[16'h2746] <= 0;
        weight_mem[16'h2747] <= 0;
        weight_mem[16'h2748] <= 0;
        weight_mem[16'h2749] <= 0;
        weight_mem[16'h274A] <= 0;
        weight_mem[16'h274B] <= 0;
        weight_mem[16'h274C] <= 0;
        weight_mem[16'h274D] <= 0;
        weight_mem[16'h274E] <= 0;
        weight_mem[16'h274F] <= 0;
        weight_mem[16'h2750] <= 0;
        weight_mem[16'h2751] <= 0;
        weight_mem[16'h2752] <= 0;
        weight_mem[16'h2753] <= 0;
        weight_mem[16'h2754] <= 0;
        weight_mem[16'h2755] <= 0;
        weight_mem[16'h2756] <= 0;
        weight_mem[16'h2757] <= 0;
        weight_mem[16'h2758] <= 0;
        weight_mem[16'h2759] <= 0;
        weight_mem[16'h275A] <= 0;
        weight_mem[16'h275B] <= 0;
        weight_mem[16'h275C] <= 0;
        weight_mem[16'h275D] <= 0;
        weight_mem[16'h275E] <= 0;
        weight_mem[16'h275F] <= 0;
        weight_mem[16'h2760] <= 0;
        weight_mem[16'h2761] <= 0;
        weight_mem[16'h2762] <= 0;
        weight_mem[16'h2763] <= 0;
        weight_mem[16'h2764] <= 0;
        weight_mem[16'h2765] <= 0;
        weight_mem[16'h2766] <= 0;
        weight_mem[16'h2767] <= 0;
        weight_mem[16'h2768] <= 0;
        weight_mem[16'h2769] <= 0;
        weight_mem[16'h276A] <= 0;
        weight_mem[16'h276B] <= 0;
        weight_mem[16'h276C] <= 0;
        weight_mem[16'h276D] <= 0;
        weight_mem[16'h276E] <= 0;
        weight_mem[16'h276F] <= 0;
        weight_mem[16'h2770] <= 0;
        weight_mem[16'h2771] <= 0;
        weight_mem[16'h2772] <= 0;
        weight_mem[16'h2773] <= 0;
        weight_mem[16'h2774] <= 0;
        weight_mem[16'h2775] <= 0;
        weight_mem[16'h2776] <= 0;
        weight_mem[16'h2777] <= 0;
        weight_mem[16'h2778] <= 0;
        weight_mem[16'h2779] <= 0;
        weight_mem[16'h277A] <= 0;
        weight_mem[16'h277B] <= 0;
        weight_mem[16'h277C] <= 0;
        weight_mem[16'h277D] <= 0;
        weight_mem[16'h277E] <= 0;
        weight_mem[16'h277F] <= 0;
        weight_mem[16'h2780] <= 0;
        weight_mem[16'h2781] <= 0;
        weight_mem[16'h2782] <= 0;
        weight_mem[16'h2783] <= 0;
        weight_mem[16'h2784] <= 0;
        weight_mem[16'h2785] <= 0;
        weight_mem[16'h2786] <= 0;
        weight_mem[16'h2787] <= 0;
        weight_mem[16'h2788] <= 0;
        weight_mem[16'h2789] <= 0;
        weight_mem[16'h278A] <= 0;
        weight_mem[16'h278B] <= 0;
        weight_mem[16'h278C] <= 0;
        weight_mem[16'h278D] <= 0;
        weight_mem[16'h278E] <= 0;
        weight_mem[16'h278F] <= 0;
        weight_mem[16'h2790] <= 0;
        weight_mem[16'h2791] <= 0;
        weight_mem[16'h2792] <= 0;
        weight_mem[16'h2793] <= 0;
        weight_mem[16'h2794] <= 0;
        weight_mem[16'h2795] <= 0;
        weight_mem[16'h2796] <= 0;
        weight_mem[16'h2797] <= 0;
        weight_mem[16'h2798] <= 0;
        weight_mem[16'h2799] <= 0;
        weight_mem[16'h279A] <= 0;
        weight_mem[16'h279B] <= 0;
        weight_mem[16'h279C] <= 0;
        weight_mem[16'h279D] <= 0;
        weight_mem[16'h279E] <= 0;
        weight_mem[16'h279F] <= 0;
        weight_mem[16'h27A0] <= 0;
        weight_mem[16'h27A1] <= 0;
        weight_mem[16'h27A2] <= 0;
        weight_mem[16'h27A3] <= 0;
        weight_mem[16'h27A4] <= 0;
        weight_mem[16'h27A5] <= 0;
        weight_mem[16'h27A6] <= 0;
        weight_mem[16'h27A7] <= 0;
        weight_mem[16'h27A8] <= 0;
        weight_mem[16'h27A9] <= 0;
        weight_mem[16'h27AA] <= 0;
        weight_mem[16'h27AB] <= 0;
        weight_mem[16'h27AC] <= 0;
        weight_mem[16'h27AD] <= 0;
        weight_mem[16'h27AE] <= 0;
        weight_mem[16'h27AF] <= 0;

        // layer 1 neuron 20
        weight_mem[16'h2800] <= 0;
        weight_mem[16'h2801] <= 0;
        weight_mem[16'h2802] <= 0;
        weight_mem[16'h2803] <= 0;
        weight_mem[16'h2804] <= 0;
        weight_mem[16'h2805] <= 0;
        weight_mem[16'h2806] <= 0;
        weight_mem[16'h2807] <= 0;
        weight_mem[16'h2808] <= 0;
        weight_mem[16'h2809] <= 0;
        weight_mem[16'h280A] <= 0;
        weight_mem[16'h280B] <= 0;
        weight_mem[16'h280C] <= 0;
        weight_mem[16'h280D] <= 0;
        weight_mem[16'h280E] <= 0;
        weight_mem[16'h280F] <= 0;
        weight_mem[16'h2810] <= 0;
        weight_mem[16'h2811] <= 0;
        weight_mem[16'h2812] <= 0;
        weight_mem[16'h2813] <= 0;
        weight_mem[16'h2814] <= 0;
        weight_mem[16'h2815] <= 0;
        weight_mem[16'h2816] <= 0;
        weight_mem[16'h2817] <= 0;
        weight_mem[16'h2818] <= 0;
        weight_mem[16'h2819] <= 0;
        weight_mem[16'h281A] <= 0;
        weight_mem[16'h281B] <= 0;
        weight_mem[16'h281C] <= 0;
        weight_mem[16'h281D] <= 0;
        weight_mem[16'h281E] <= 0;
        weight_mem[16'h281F] <= 0;
        weight_mem[16'h2820] <= 0;
        weight_mem[16'h2821] <= 0;
        weight_mem[16'h2822] <= 0;
        weight_mem[16'h2823] <= 0;
        weight_mem[16'h2824] <= 0;
        weight_mem[16'h2825] <= 0;
        weight_mem[16'h2826] <= 0;
        weight_mem[16'h2827] <= 0;
        weight_mem[16'h2828] <= 0;
        weight_mem[16'h2829] <= 0;
        weight_mem[16'h282A] <= 0;
        weight_mem[16'h282B] <= 0;
        weight_mem[16'h282C] <= 0;
        weight_mem[16'h282D] <= 0;
        weight_mem[16'h282E] <= 0;
        weight_mem[16'h282F] <= 0;
        weight_mem[16'h2830] <= 0;
        weight_mem[16'h2831] <= 0;
        weight_mem[16'h2832] <= 0;
        weight_mem[16'h2833] <= 0;
        weight_mem[16'h2834] <= 0;
        weight_mem[16'h2835] <= 0;
        weight_mem[16'h2836] <= 0;
        weight_mem[16'h2837] <= 0;
        weight_mem[16'h2838] <= 0;
        weight_mem[16'h2839] <= 0;
        weight_mem[16'h283A] <= 0;
        weight_mem[16'h283B] <= 0;
        weight_mem[16'h283C] <= 0;
        weight_mem[16'h283D] <= 0;
        weight_mem[16'h283E] <= 0;
        weight_mem[16'h283F] <= 0;
        weight_mem[16'h2840] <= 0;
        weight_mem[16'h2841] <= 0;
        weight_mem[16'h2842] <= 0;
        weight_mem[16'h2843] <= 0;
        weight_mem[16'h2844] <= 0;
        weight_mem[16'h2845] <= 0;
        weight_mem[16'h2846] <= 0;
        weight_mem[16'h2847] <= 0;
        weight_mem[16'h2848] <= 0;
        weight_mem[16'h2849] <= 0;
        weight_mem[16'h284A] <= 0;
        weight_mem[16'h284B] <= 0;
        weight_mem[16'h284C] <= 0;
        weight_mem[16'h284D] <= 0;
        weight_mem[16'h284E] <= 0;
        weight_mem[16'h284F] <= 0;
        weight_mem[16'h2850] <= 0;
        weight_mem[16'h2851] <= 0;
        weight_mem[16'h2852] <= 0;
        weight_mem[16'h2853] <= 0;
        weight_mem[16'h2854] <= 0;
        weight_mem[16'h2855] <= 0;
        weight_mem[16'h2856] <= 0;
        weight_mem[16'h2857] <= 0;
        weight_mem[16'h2858] <= 0;
        weight_mem[16'h2859] <= 0;
        weight_mem[16'h285A] <= 0;
        weight_mem[16'h285B] <= 0;
        weight_mem[16'h285C] <= 0;
        weight_mem[16'h285D] <= 0;
        weight_mem[16'h285E] <= 0;
        weight_mem[16'h285F] <= 0;
        weight_mem[16'h2860] <= 0;
        weight_mem[16'h2861] <= 0;
        weight_mem[16'h2862] <= 0;
        weight_mem[16'h2863] <= 0;
        weight_mem[16'h2864] <= 0;
        weight_mem[16'h2865] <= 0;
        weight_mem[16'h2866] <= 0;
        weight_mem[16'h2867] <= 0;
        weight_mem[16'h2868] <= 0;
        weight_mem[16'h2869] <= 0;
        weight_mem[16'h286A] <= 0;
        weight_mem[16'h286B] <= 0;
        weight_mem[16'h286C] <= 0;
        weight_mem[16'h286D] <= 0;
        weight_mem[16'h286E] <= 0;
        weight_mem[16'h286F] <= 0;
        weight_mem[16'h2870] <= 0;
        weight_mem[16'h2871] <= 0;
        weight_mem[16'h2872] <= 0;
        weight_mem[16'h2873] <= 0;
        weight_mem[16'h2874] <= 0;
        weight_mem[16'h2875] <= 0;
        weight_mem[16'h2876] <= 0;
        weight_mem[16'h2877] <= 0;
        weight_mem[16'h2878] <= 0;
        weight_mem[16'h2879] <= 0;
        weight_mem[16'h287A] <= 0;
        weight_mem[16'h287B] <= 0;
        weight_mem[16'h287C] <= 0;
        weight_mem[16'h287D] <= 0;
        weight_mem[16'h287E] <= 0;
        weight_mem[16'h287F] <= 0;
        weight_mem[16'h2880] <= 0;
        weight_mem[16'h2881] <= 0;
        weight_mem[16'h2882] <= 0;
        weight_mem[16'h2883] <= 0;
        weight_mem[16'h2884] <= 0;
        weight_mem[16'h2885] <= 0;
        weight_mem[16'h2886] <= 0;
        weight_mem[16'h2887] <= 0;
        weight_mem[16'h2888] <= 0;
        weight_mem[16'h2889] <= 0;
        weight_mem[16'h288A] <= 0;
        weight_mem[16'h288B] <= 0;
        weight_mem[16'h288C] <= 0;
        weight_mem[16'h288D] <= 0;
        weight_mem[16'h288E] <= 0;
        weight_mem[16'h288F] <= 0;
        weight_mem[16'h2890] <= 0;
        weight_mem[16'h2891] <= 0;
        weight_mem[16'h2892] <= 0;
        weight_mem[16'h2893] <= 0;
        weight_mem[16'h2894] <= 0;
        weight_mem[16'h2895] <= 0;
        weight_mem[16'h2896] <= 0;
        weight_mem[16'h2897] <= 0;
        weight_mem[16'h2898] <= 0;
        weight_mem[16'h2899] <= 0;
        weight_mem[16'h289A] <= 0;
        weight_mem[16'h289B] <= 0;
        weight_mem[16'h289C] <= 0;
        weight_mem[16'h289D] <= 0;
        weight_mem[16'h289E] <= 0;
        weight_mem[16'h289F] <= 0;
        weight_mem[16'h28A0] <= 0;
        weight_mem[16'h28A1] <= 0;
        weight_mem[16'h28A2] <= 0;
        weight_mem[16'h28A3] <= 0;
        weight_mem[16'h28A4] <= 0;
        weight_mem[16'h28A5] <= 0;
        weight_mem[16'h28A6] <= 0;
        weight_mem[16'h28A7] <= 0;
        weight_mem[16'h28A8] <= 0;
        weight_mem[16'h28A9] <= 0;
        weight_mem[16'h28AA] <= 0;
        weight_mem[16'h28AB] <= 0;
        weight_mem[16'h28AC] <= 0;
        weight_mem[16'h28AD] <= 0;
        weight_mem[16'h28AE] <= 0;
        weight_mem[16'h28AF] <= 0;
        weight_mem[16'h28B0] <= 0;
        weight_mem[16'h28B1] <= 0;
        weight_mem[16'h28B2] <= 0;
        weight_mem[16'h28B3] <= 0;
        weight_mem[16'h28B4] <= 0;
        weight_mem[16'h28B5] <= 0;
        weight_mem[16'h28B6] <= 0;
        weight_mem[16'h28B7] <= 0;
        weight_mem[16'h28B8] <= 0;
        weight_mem[16'h28B9] <= 0;
        weight_mem[16'h28BA] <= 0;
        weight_mem[16'h28BB] <= 0;
        weight_mem[16'h28BC] <= 0;
        weight_mem[16'h28BD] <= 0;
        weight_mem[16'h28BE] <= 0;
        weight_mem[16'h28BF] <= 0;
        weight_mem[16'h28C0] <= 0;
        weight_mem[16'h28C1] <= 0;
        weight_mem[16'h28C2] <= 0;
        weight_mem[16'h28C3] <= 0;
        weight_mem[16'h28C4] <= 0;
        weight_mem[16'h28C5] <= 0;
        weight_mem[16'h28C6] <= 0;
        weight_mem[16'h28C7] <= 0;
        weight_mem[16'h28C8] <= 0;
        weight_mem[16'h28C9] <= 0;
        weight_mem[16'h28CA] <= 0;
        weight_mem[16'h28CB] <= 0;
        weight_mem[16'h28CC] <= 0;
        weight_mem[16'h28CD] <= 0;
        weight_mem[16'h28CE] <= 0;
        weight_mem[16'h28CF] <= 0;
        weight_mem[16'h28D0] <= 0;
        weight_mem[16'h28D1] <= 0;
        weight_mem[16'h28D2] <= 0;
        weight_mem[16'h28D3] <= 0;
        weight_mem[16'h28D4] <= 0;
        weight_mem[16'h28D5] <= 0;
        weight_mem[16'h28D6] <= 0;
        weight_mem[16'h28D7] <= 0;
        weight_mem[16'h28D8] <= 0;
        weight_mem[16'h28D9] <= 0;
        weight_mem[16'h28DA] <= 0;
        weight_mem[16'h28DB] <= 0;
        weight_mem[16'h28DC] <= 0;
        weight_mem[16'h28DD] <= 0;
        weight_mem[16'h28DE] <= 0;
        weight_mem[16'h28DF] <= 0;
        weight_mem[16'h28E0] <= 0;
        weight_mem[16'h28E1] <= 0;
        weight_mem[16'h28E2] <= 0;
        weight_mem[16'h28E3] <= 0;
        weight_mem[16'h28E4] <= 0;
        weight_mem[16'h28E5] <= 0;
        weight_mem[16'h28E6] <= 0;
        weight_mem[16'h28E7] <= 0;
        weight_mem[16'h28E8] <= 0;
        weight_mem[16'h28E9] <= 0;
        weight_mem[16'h28EA] <= 0;
        weight_mem[16'h28EB] <= 0;
        weight_mem[16'h28EC] <= 0;
        weight_mem[16'h28ED] <= 0;
        weight_mem[16'h28EE] <= 0;
        weight_mem[16'h28EF] <= 0;
        weight_mem[16'h28F0] <= 0;
        weight_mem[16'h28F1] <= 0;
        weight_mem[16'h28F2] <= 0;
        weight_mem[16'h28F3] <= 0;
        weight_mem[16'h28F4] <= 0;
        weight_mem[16'h28F5] <= 0;
        weight_mem[16'h28F6] <= 0;
        weight_mem[16'h28F7] <= 0;
        weight_mem[16'h28F8] <= 0;
        weight_mem[16'h28F9] <= 0;
        weight_mem[16'h28FA] <= 0;
        weight_mem[16'h28FB] <= 0;
        weight_mem[16'h28FC] <= 0;
        weight_mem[16'h28FD] <= 0;
        weight_mem[16'h28FE] <= 0;
        weight_mem[16'h28FF] <= 0;
        weight_mem[16'h2900] <= 0;
        weight_mem[16'h2901] <= 0;
        weight_mem[16'h2902] <= 0;
        weight_mem[16'h2903] <= 0;
        weight_mem[16'h2904] <= 0;
        weight_mem[16'h2905] <= 0;
        weight_mem[16'h2906] <= 0;
        weight_mem[16'h2907] <= 0;
        weight_mem[16'h2908] <= 0;
        weight_mem[16'h2909] <= 0;
        weight_mem[16'h290A] <= 0;
        weight_mem[16'h290B] <= 0;
        weight_mem[16'h290C] <= 0;
        weight_mem[16'h290D] <= 0;
        weight_mem[16'h290E] <= 0;
        weight_mem[16'h290F] <= 0;
        weight_mem[16'h2910] <= 0;
        weight_mem[16'h2911] <= 0;
        weight_mem[16'h2912] <= 0;
        weight_mem[16'h2913] <= 0;
        weight_mem[16'h2914] <= 0;
        weight_mem[16'h2915] <= 0;
        weight_mem[16'h2916] <= 0;
        weight_mem[16'h2917] <= 0;
        weight_mem[16'h2918] <= 0;
        weight_mem[16'h2919] <= 0;
        weight_mem[16'h291A] <= 0;
        weight_mem[16'h291B] <= 0;
        weight_mem[16'h291C] <= 0;
        weight_mem[16'h291D] <= 0;
        weight_mem[16'h291E] <= 0;
        weight_mem[16'h291F] <= 0;
        weight_mem[16'h2920] <= 0;
        weight_mem[16'h2921] <= 0;
        weight_mem[16'h2922] <= 0;
        weight_mem[16'h2923] <= 0;
        weight_mem[16'h2924] <= 0;
        weight_mem[16'h2925] <= 0;
        weight_mem[16'h2926] <= 0;
        weight_mem[16'h2927] <= 0;
        weight_mem[16'h2928] <= 0;
        weight_mem[16'h2929] <= 0;
        weight_mem[16'h292A] <= 0;
        weight_mem[16'h292B] <= 0;
        weight_mem[16'h292C] <= 0;
        weight_mem[16'h292D] <= 0;
        weight_mem[16'h292E] <= 0;
        weight_mem[16'h292F] <= 0;
        weight_mem[16'h2930] <= 0;
        weight_mem[16'h2931] <= 0;
        weight_mem[16'h2932] <= 0;
        weight_mem[16'h2933] <= 0;
        weight_mem[16'h2934] <= 0;
        weight_mem[16'h2935] <= 0;
        weight_mem[16'h2936] <= 0;
        weight_mem[16'h2937] <= 0;
        weight_mem[16'h2938] <= 0;
        weight_mem[16'h2939] <= 0;
        weight_mem[16'h293A] <= 0;
        weight_mem[16'h293B] <= 0;
        weight_mem[16'h293C] <= 0;
        weight_mem[16'h293D] <= 0;
        weight_mem[16'h293E] <= 0;
        weight_mem[16'h293F] <= 0;
        weight_mem[16'h2940] <= 0;
        weight_mem[16'h2941] <= 0;
        weight_mem[16'h2942] <= 0;
        weight_mem[16'h2943] <= 0;
        weight_mem[16'h2944] <= 0;
        weight_mem[16'h2945] <= 0;
        weight_mem[16'h2946] <= 0;
        weight_mem[16'h2947] <= 0;
        weight_mem[16'h2948] <= 0;
        weight_mem[16'h2949] <= 0;
        weight_mem[16'h294A] <= 0;
        weight_mem[16'h294B] <= 0;
        weight_mem[16'h294C] <= 0;
        weight_mem[16'h294D] <= 0;
        weight_mem[16'h294E] <= 0;
        weight_mem[16'h294F] <= 0;
        weight_mem[16'h2950] <= 0;
        weight_mem[16'h2951] <= 0;
        weight_mem[16'h2952] <= 0;
        weight_mem[16'h2953] <= 0;
        weight_mem[16'h2954] <= 0;
        weight_mem[16'h2955] <= 0;
        weight_mem[16'h2956] <= 0;
        weight_mem[16'h2957] <= 0;
        weight_mem[16'h2958] <= 0;
        weight_mem[16'h2959] <= 0;
        weight_mem[16'h295A] <= 0;
        weight_mem[16'h295B] <= 0;
        weight_mem[16'h295C] <= 0;
        weight_mem[16'h295D] <= 0;
        weight_mem[16'h295E] <= 0;
        weight_mem[16'h295F] <= 0;
        weight_mem[16'h2960] <= 0;
        weight_mem[16'h2961] <= 0;
        weight_mem[16'h2962] <= 0;
        weight_mem[16'h2963] <= 0;
        weight_mem[16'h2964] <= 0;
        weight_mem[16'h2965] <= 0;
        weight_mem[16'h2966] <= 0;
        weight_mem[16'h2967] <= 0;
        weight_mem[16'h2968] <= 0;
        weight_mem[16'h2969] <= 0;
        weight_mem[16'h296A] <= 0;
        weight_mem[16'h296B] <= 0;
        weight_mem[16'h296C] <= 0;
        weight_mem[16'h296D] <= 0;
        weight_mem[16'h296E] <= 0;
        weight_mem[16'h296F] <= 0;
        weight_mem[16'h2970] <= 0;
        weight_mem[16'h2971] <= 0;
        weight_mem[16'h2972] <= 0;
        weight_mem[16'h2973] <= 0;
        weight_mem[16'h2974] <= 0;
        weight_mem[16'h2975] <= 0;
        weight_mem[16'h2976] <= 0;
        weight_mem[16'h2977] <= 0;
        weight_mem[16'h2978] <= 0;
        weight_mem[16'h2979] <= 0;
        weight_mem[16'h297A] <= 0;
        weight_mem[16'h297B] <= 0;
        weight_mem[16'h297C] <= 0;
        weight_mem[16'h297D] <= 0;
        weight_mem[16'h297E] <= 0;
        weight_mem[16'h297F] <= 0;
        weight_mem[16'h2980] <= 0;
        weight_mem[16'h2981] <= 0;
        weight_mem[16'h2982] <= 0;
        weight_mem[16'h2983] <= 0;
        weight_mem[16'h2984] <= 0;
        weight_mem[16'h2985] <= 0;
        weight_mem[16'h2986] <= 0;
        weight_mem[16'h2987] <= 0;
        weight_mem[16'h2988] <= 0;
        weight_mem[16'h2989] <= 0;
        weight_mem[16'h298A] <= 0;
        weight_mem[16'h298B] <= 0;
        weight_mem[16'h298C] <= 0;
        weight_mem[16'h298D] <= 0;
        weight_mem[16'h298E] <= 0;
        weight_mem[16'h298F] <= 0;
        weight_mem[16'h2990] <= 0;
        weight_mem[16'h2991] <= 0;
        weight_mem[16'h2992] <= 0;
        weight_mem[16'h2993] <= 0;
        weight_mem[16'h2994] <= 0;
        weight_mem[16'h2995] <= 0;
        weight_mem[16'h2996] <= 0;
        weight_mem[16'h2997] <= 0;
        weight_mem[16'h2998] <= 0;
        weight_mem[16'h2999] <= 0;
        weight_mem[16'h299A] <= 0;
        weight_mem[16'h299B] <= 0;
        weight_mem[16'h299C] <= 0;
        weight_mem[16'h299D] <= 0;
        weight_mem[16'h299E] <= 0;
        weight_mem[16'h299F] <= 0;
        weight_mem[16'h29A0] <= 0;
        weight_mem[16'h29A1] <= 0;
        weight_mem[16'h29A2] <= 0;
        weight_mem[16'h29A3] <= 0;
        weight_mem[16'h29A4] <= 0;
        weight_mem[16'h29A5] <= 0;
        weight_mem[16'h29A6] <= 0;
        weight_mem[16'h29A7] <= 0;
        weight_mem[16'h29A8] <= 0;
        weight_mem[16'h29A9] <= 0;
        weight_mem[16'h29AA] <= 0;
        weight_mem[16'h29AB] <= 0;
        weight_mem[16'h29AC] <= 0;
        weight_mem[16'h29AD] <= 0;
        weight_mem[16'h29AE] <= 0;
        weight_mem[16'h29AF] <= 0;

        // layer 1 neuron 21
        weight_mem[16'h2A00] <= 0;
        weight_mem[16'h2A01] <= 0;
        weight_mem[16'h2A02] <= 0;
        weight_mem[16'h2A03] <= 0;
        weight_mem[16'h2A04] <= 0;
        weight_mem[16'h2A05] <= 0;
        weight_mem[16'h2A06] <= 0;
        weight_mem[16'h2A07] <= 0;
        weight_mem[16'h2A08] <= 0;
        weight_mem[16'h2A09] <= 0;
        weight_mem[16'h2A0A] <= 0;
        weight_mem[16'h2A0B] <= 0;
        weight_mem[16'h2A0C] <= 0;
        weight_mem[16'h2A0D] <= 0;
        weight_mem[16'h2A0E] <= 0;
        weight_mem[16'h2A0F] <= 0;
        weight_mem[16'h2A10] <= 0;
        weight_mem[16'h2A11] <= 0;
        weight_mem[16'h2A12] <= 0;
        weight_mem[16'h2A13] <= 0;
        weight_mem[16'h2A14] <= 0;
        weight_mem[16'h2A15] <= 0;
        weight_mem[16'h2A16] <= 0;
        weight_mem[16'h2A17] <= 0;
        weight_mem[16'h2A18] <= 0;
        weight_mem[16'h2A19] <= 0;
        weight_mem[16'h2A1A] <= 0;
        weight_mem[16'h2A1B] <= 0;
        weight_mem[16'h2A1C] <= 0;
        weight_mem[16'h2A1D] <= 0;
        weight_mem[16'h2A1E] <= 0;
        weight_mem[16'h2A1F] <= 0;
        weight_mem[16'h2A20] <= 0;
        weight_mem[16'h2A21] <= 0;
        weight_mem[16'h2A22] <= 0;
        weight_mem[16'h2A23] <= 0;
        weight_mem[16'h2A24] <= 0;
        weight_mem[16'h2A25] <= 0;
        weight_mem[16'h2A26] <= 0;
        weight_mem[16'h2A27] <= 0;
        weight_mem[16'h2A28] <= 0;
        weight_mem[16'h2A29] <= 0;
        weight_mem[16'h2A2A] <= 0;
        weight_mem[16'h2A2B] <= 0;
        weight_mem[16'h2A2C] <= 0;
        weight_mem[16'h2A2D] <= 0;
        weight_mem[16'h2A2E] <= 0;
        weight_mem[16'h2A2F] <= 0;
        weight_mem[16'h2A30] <= 0;
        weight_mem[16'h2A31] <= 0;
        weight_mem[16'h2A32] <= 0;
        weight_mem[16'h2A33] <= 0;
        weight_mem[16'h2A34] <= 0;
        weight_mem[16'h2A35] <= 0;
        weight_mem[16'h2A36] <= 0;
        weight_mem[16'h2A37] <= 0;
        weight_mem[16'h2A38] <= 0;
        weight_mem[16'h2A39] <= 0;
        weight_mem[16'h2A3A] <= 0;
        weight_mem[16'h2A3B] <= 0;
        weight_mem[16'h2A3C] <= 0;
        weight_mem[16'h2A3D] <= 0;
        weight_mem[16'h2A3E] <= 0;
        weight_mem[16'h2A3F] <= 0;
        weight_mem[16'h2A40] <= 0;
        weight_mem[16'h2A41] <= 0;
        weight_mem[16'h2A42] <= 0;
        weight_mem[16'h2A43] <= 0;
        weight_mem[16'h2A44] <= 0;
        weight_mem[16'h2A45] <= 0;
        weight_mem[16'h2A46] <= 0;
        weight_mem[16'h2A47] <= 0;
        weight_mem[16'h2A48] <= 0;
        weight_mem[16'h2A49] <= 0;
        weight_mem[16'h2A4A] <= 0;
        weight_mem[16'h2A4B] <= 0;
        weight_mem[16'h2A4C] <= 0;
        weight_mem[16'h2A4D] <= 0;
        weight_mem[16'h2A4E] <= 0;
        weight_mem[16'h2A4F] <= 0;
        weight_mem[16'h2A50] <= 0;
        weight_mem[16'h2A51] <= 0;
        weight_mem[16'h2A52] <= 0;
        weight_mem[16'h2A53] <= 0;
        weight_mem[16'h2A54] <= 0;
        weight_mem[16'h2A55] <= 0;
        weight_mem[16'h2A56] <= 0;
        weight_mem[16'h2A57] <= 0;
        weight_mem[16'h2A58] <= 0;
        weight_mem[16'h2A59] <= 0;
        weight_mem[16'h2A5A] <= 0;
        weight_mem[16'h2A5B] <= 0;
        weight_mem[16'h2A5C] <= 0;
        weight_mem[16'h2A5D] <= 0;
        weight_mem[16'h2A5E] <= 0;
        weight_mem[16'h2A5F] <= 0;
        weight_mem[16'h2A60] <= 0;
        weight_mem[16'h2A61] <= 0;
        weight_mem[16'h2A62] <= 0;
        weight_mem[16'h2A63] <= 0;
        weight_mem[16'h2A64] <= 0;
        weight_mem[16'h2A65] <= 0;
        weight_mem[16'h2A66] <= 0;
        weight_mem[16'h2A67] <= 0;
        weight_mem[16'h2A68] <= 0;
        weight_mem[16'h2A69] <= 0;
        weight_mem[16'h2A6A] <= 0;
        weight_mem[16'h2A6B] <= 0;
        weight_mem[16'h2A6C] <= 0;
        weight_mem[16'h2A6D] <= 0;
        weight_mem[16'h2A6E] <= 0;
        weight_mem[16'h2A6F] <= 0;
        weight_mem[16'h2A70] <= 0;
        weight_mem[16'h2A71] <= 0;
        weight_mem[16'h2A72] <= 0;
        weight_mem[16'h2A73] <= 0;
        weight_mem[16'h2A74] <= 0;
        weight_mem[16'h2A75] <= 0;
        weight_mem[16'h2A76] <= 0;
        weight_mem[16'h2A77] <= 0;
        weight_mem[16'h2A78] <= 0;
        weight_mem[16'h2A79] <= 0;
        weight_mem[16'h2A7A] <= 0;
        weight_mem[16'h2A7B] <= 0;
        weight_mem[16'h2A7C] <= 0;
        weight_mem[16'h2A7D] <= 0;
        weight_mem[16'h2A7E] <= 0;
        weight_mem[16'h2A7F] <= 0;
        weight_mem[16'h2A80] <= 0;
        weight_mem[16'h2A81] <= 0;
        weight_mem[16'h2A82] <= 0;
        weight_mem[16'h2A83] <= 0;
        weight_mem[16'h2A84] <= 0;
        weight_mem[16'h2A85] <= 0;
        weight_mem[16'h2A86] <= 0;
        weight_mem[16'h2A87] <= 0;
        weight_mem[16'h2A88] <= 0;
        weight_mem[16'h2A89] <= 0;
        weight_mem[16'h2A8A] <= 0;
        weight_mem[16'h2A8B] <= 0;
        weight_mem[16'h2A8C] <= 0;
        weight_mem[16'h2A8D] <= 0;
        weight_mem[16'h2A8E] <= 0;
        weight_mem[16'h2A8F] <= 0;
        weight_mem[16'h2A90] <= 0;
        weight_mem[16'h2A91] <= 0;
        weight_mem[16'h2A92] <= 0;
        weight_mem[16'h2A93] <= 0;
        weight_mem[16'h2A94] <= 0;
        weight_mem[16'h2A95] <= 0;
        weight_mem[16'h2A96] <= 0;
        weight_mem[16'h2A97] <= 0;
        weight_mem[16'h2A98] <= 0;
        weight_mem[16'h2A99] <= 0;
        weight_mem[16'h2A9A] <= 0;
        weight_mem[16'h2A9B] <= 0;
        weight_mem[16'h2A9C] <= 0;
        weight_mem[16'h2A9D] <= 0;
        weight_mem[16'h2A9E] <= 0;
        weight_mem[16'h2A9F] <= 0;
        weight_mem[16'h2AA0] <= 0;
        weight_mem[16'h2AA1] <= 0;
        weight_mem[16'h2AA2] <= 0;
        weight_mem[16'h2AA3] <= 0;
        weight_mem[16'h2AA4] <= 0;
        weight_mem[16'h2AA5] <= 0;
        weight_mem[16'h2AA6] <= 0;
        weight_mem[16'h2AA7] <= 0;
        weight_mem[16'h2AA8] <= 0;
        weight_mem[16'h2AA9] <= 0;
        weight_mem[16'h2AAA] <= 0;
        weight_mem[16'h2AAB] <= 0;
        weight_mem[16'h2AAC] <= 0;
        weight_mem[16'h2AAD] <= 0;
        weight_mem[16'h2AAE] <= 0;
        weight_mem[16'h2AAF] <= 0;
        weight_mem[16'h2AB0] <= 0;
        weight_mem[16'h2AB1] <= 0;
        weight_mem[16'h2AB2] <= 0;
        weight_mem[16'h2AB3] <= 0;
        weight_mem[16'h2AB4] <= 0;
        weight_mem[16'h2AB5] <= 0;
        weight_mem[16'h2AB6] <= 0;
        weight_mem[16'h2AB7] <= 0;
        weight_mem[16'h2AB8] <= 0;
        weight_mem[16'h2AB9] <= 0;
        weight_mem[16'h2ABA] <= 0;
        weight_mem[16'h2ABB] <= 0;
        weight_mem[16'h2ABC] <= 0;
        weight_mem[16'h2ABD] <= 0;
        weight_mem[16'h2ABE] <= 0;
        weight_mem[16'h2ABF] <= 0;
        weight_mem[16'h2AC0] <= 0;
        weight_mem[16'h2AC1] <= 0;
        weight_mem[16'h2AC2] <= 0;
        weight_mem[16'h2AC3] <= 0;
        weight_mem[16'h2AC4] <= 0;
        weight_mem[16'h2AC5] <= 0;
        weight_mem[16'h2AC6] <= 0;
        weight_mem[16'h2AC7] <= 0;
        weight_mem[16'h2AC8] <= 0;
        weight_mem[16'h2AC9] <= 0;
        weight_mem[16'h2ACA] <= 0;
        weight_mem[16'h2ACB] <= 0;
        weight_mem[16'h2ACC] <= 0;
        weight_mem[16'h2ACD] <= 0;
        weight_mem[16'h2ACE] <= 0;
        weight_mem[16'h2ACF] <= 0;
        weight_mem[16'h2AD0] <= 0;
        weight_mem[16'h2AD1] <= 0;
        weight_mem[16'h2AD2] <= 0;
        weight_mem[16'h2AD3] <= 0;
        weight_mem[16'h2AD4] <= 0;
        weight_mem[16'h2AD5] <= 0;
        weight_mem[16'h2AD6] <= 0;
        weight_mem[16'h2AD7] <= 0;
        weight_mem[16'h2AD8] <= 0;
        weight_mem[16'h2AD9] <= 0;
        weight_mem[16'h2ADA] <= 0;
        weight_mem[16'h2ADB] <= 0;
        weight_mem[16'h2ADC] <= 0;
        weight_mem[16'h2ADD] <= 0;
        weight_mem[16'h2ADE] <= 0;
        weight_mem[16'h2ADF] <= 0;
        weight_mem[16'h2AE0] <= 0;
        weight_mem[16'h2AE1] <= 0;
        weight_mem[16'h2AE2] <= 0;
        weight_mem[16'h2AE3] <= 0;
        weight_mem[16'h2AE4] <= 0;
        weight_mem[16'h2AE5] <= 0;
        weight_mem[16'h2AE6] <= 0;
        weight_mem[16'h2AE7] <= 0;
        weight_mem[16'h2AE8] <= 0;
        weight_mem[16'h2AE9] <= 0;
        weight_mem[16'h2AEA] <= 0;
        weight_mem[16'h2AEB] <= 0;
        weight_mem[16'h2AEC] <= 0;
        weight_mem[16'h2AED] <= 0;
        weight_mem[16'h2AEE] <= 0;
        weight_mem[16'h2AEF] <= 0;
        weight_mem[16'h2AF0] <= 0;
        weight_mem[16'h2AF1] <= 0;
        weight_mem[16'h2AF2] <= 0;
        weight_mem[16'h2AF3] <= 0;
        weight_mem[16'h2AF4] <= 0;
        weight_mem[16'h2AF5] <= 0;
        weight_mem[16'h2AF6] <= 0;
        weight_mem[16'h2AF7] <= 0;
        weight_mem[16'h2AF8] <= 0;
        weight_mem[16'h2AF9] <= 0;
        weight_mem[16'h2AFA] <= 0;
        weight_mem[16'h2AFB] <= 0;
        weight_mem[16'h2AFC] <= 0;
        weight_mem[16'h2AFD] <= 0;
        weight_mem[16'h2AFE] <= 0;
        weight_mem[16'h2AFF] <= 0;
        weight_mem[16'h2B00] <= 0;
        weight_mem[16'h2B01] <= 0;
        weight_mem[16'h2B02] <= 0;
        weight_mem[16'h2B03] <= 0;
        weight_mem[16'h2B04] <= 0;
        weight_mem[16'h2B05] <= 0;
        weight_mem[16'h2B06] <= 0;
        weight_mem[16'h2B07] <= 0;
        weight_mem[16'h2B08] <= 0;
        weight_mem[16'h2B09] <= 0;
        weight_mem[16'h2B0A] <= 0;
        weight_mem[16'h2B0B] <= 0;
        weight_mem[16'h2B0C] <= 0;
        weight_mem[16'h2B0D] <= 0;
        weight_mem[16'h2B0E] <= 0;
        weight_mem[16'h2B0F] <= 0;
        weight_mem[16'h2B10] <= 0;
        weight_mem[16'h2B11] <= 0;
        weight_mem[16'h2B12] <= 0;
        weight_mem[16'h2B13] <= 0;
        weight_mem[16'h2B14] <= 0;
        weight_mem[16'h2B15] <= 0;
        weight_mem[16'h2B16] <= 0;
        weight_mem[16'h2B17] <= 0;
        weight_mem[16'h2B18] <= 0;
        weight_mem[16'h2B19] <= 0;
        weight_mem[16'h2B1A] <= 0;
        weight_mem[16'h2B1B] <= 0;
        weight_mem[16'h2B1C] <= 0;
        weight_mem[16'h2B1D] <= 0;
        weight_mem[16'h2B1E] <= 0;
        weight_mem[16'h2B1F] <= 0;
        weight_mem[16'h2B20] <= 0;
        weight_mem[16'h2B21] <= 0;
        weight_mem[16'h2B22] <= 0;
        weight_mem[16'h2B23] <= 0;
        weight_mem[16'h2B24] <= 0;
        weight_mem[16'h2B25] <= 0;
        weight_mem[16'h2B26] <= 0;
        weight_mem[16'h2B27] <= 0;
        weight_mem[16'h2B28] <= 0;
        weight_mem[16'h2B29] <= 0;
        weight_mem[16'h2B2A] <= 0;
        weight_mem[16'h2B2B] <= 0;
        weight_mem[16'h2B2C] <= 0;
        weight_mem[16'h2B2D] <= 0;
        weight_mem[16'h2B2E] <= 0;
        weight_mem[16'h2B2F] <= 0;
        weight_mem[16'h2B30] <= 0;
        weight_mem[16'h2B31] <= 0;
        weight_mem[16'h2B32] <= 0;
        weight_mem[16'h2B33] <= 0;
        weight_mem[16'h2B34] <= 0;
        weight_mem[16'h2B35] <= 0;
        weight_mem[16'h2B36] <= 0;
        weight_mem[16'h2B37] <= 0;
        weight_mem[16'h2B38] <= 0;
        weight_mem[16'h2B39] <= 0;
        weight_mem[16'h2B3A] <= 0;
        weight_mem[16'h2B3B] <= 0;
        weight_mem[16'h2B3C] <= 0;
        weight_mem[16'h2B3D] <= 0;
        weight_mem[16'h2B3E] <= 0;
        weight_mem[16'h2B3F] <= 0;
        weight_mem[16'h2B40] <= 0;
        weight_mem[16'h2B41] <= 0;
        weight_mem[16'h2B42] <= 0;
        weight_mem[16'h2B43] <= 0;
        weight_mem[16'h2B44] <= 0;
        weight_mem[16'h2B45] <= 0;
        weight_mem[16'h2B46] <= 0;
        weight_mem[16'h2B47] <= 0;
        weight_mem[16'h2B48] <= 0;
        weight_mem[16'h2B49] <= 0;
        weight_mem[16'h2B4A] <= 0;
        weight_mem[16'h2B4B] <= 0;
        weight_mem[16'h2B4C] <= 0;
        weight_mem[16'h2B4D] <= 0;
        weight_mem[16'h2B4E] <= 0;
        weight_mem[16'h2B4F] <= 0;
        weight_mem[16'h2B50] <= 0;
        weight_mem[16'h2B51] <= 0;
        weight_mem[16'h2B52] <= 0;
        weight_mem[16'h2B53] <= 0;
        weight_mem[16'h2B54] <= 0;
        weight_mem[16'h2B55] <= 0;
        weight_mem[16'h2B56] <= 0;
        weight_mem[16'h2B57] <= 0;
        weight_mem[16'h2B58] <= 0;
        weight_mem[16'h2B59] <= 0;
        weight_mem[16'h2B5A] <= 0;
        weight_mem[16'h2B5B] <= 0;
        weight_mem[16'h2B5C] <= 0;
        weight_mem[16'h2B5D] <= 0;
        weight_mem[16'h2B5E] <= 0;
        weight_mem[16'h2B5F] <= 0;
        weight_mem[16'h2B60] <= 0;
        weight_mem[16'h2B61] <= 0;
        weight_mem[16'h2B62] <= 0;
        weight_mem[16'h2B63] <= 0;
        weight_mem[16'h2B64] <= 0;
        weight_mem[16'h2B65] <= 0;
        weight_mem[16'h2B66] <= 0;
        weight_mem[16'h2B67] <= 0;
        weight_mem[16'h2B68] <= 0;
        weight_mem[16'h2B69] <= 0;
        weight_mem[16'h2B6A] <= 0;
        weight_mem[16'h2B6B] <= 0;
        weight_mem[16'h2B6C] <= 0;
        weight_mem[16'h2B6D] <= 0;
        weight_mem[16'h2B6E] <= 0;
        weight_mem[16'h2B6F] <= 0;
        weight_mem[16'h2B70] <= 0;
        weight_mem[16'h2B71] <= 0;
        weight_mem[16'h2B72] <= 0;
        weight_mem[16'h2B73] <= 0;
        weight_mem[16'h2B74] <= 0;
        weight_mem[16'h2B75] <= 0;
        weight_mem[16'h2B76] <= 0;
        weight_mem[16'h2B77] <= 0;
        weight_mem[16'h2B78] <= 0;
        weight_mem[16'h2B79] <= 0;
        weight_mem[16'h2B7A] <= 0;
        weight_mem[16'h2B7B] <= 0;
        weight_mem[16'h2B7C] <= 0;
        weight_mem[16'h2B7D] <= 0;
        weight_mem[16'h2B7E] <= 0;
        weight_mem[16'h2B7F] <= 0;
        weight_mem[16'h2B80] <= 0;
        weight_mem[16'h2B81] <= 0;
        weight_mem[16'h2B82] <= 0;
        weight_mem[16'h2B83] <= 0;
        weight_mem[16'h2B84] <= 0;
        weight_mem[16'h2B85] <= 0;
        weight_mem[16'h2B86] <= 0;
        weight_mem[16'h2B87] <= 0;
        weight_mem[16'h2B88] <= 0;
        weight_mem[16'h2B89] <= 0;
        weight_mem[16'h2B8A] <= 0;
        weight_mem[16'h2B8B] <= 0;
        weight_mem[16'h2B8C] <= 0;
        weight_mem[16'h2B8D] <= 0;
        weight_mem[16'h2B8E] <= 0;
        weight_mem[16'h2B8F] <= 0;
        weight_mem[16'h2B90] <= 0;
        weight_mem[16'h2B91] <= 0;
        weight_mem[16'h2B92] <= 0;
        weight_mem[16'h2B93] <= 0;
        weight_mem[16'h2B94] <= 0;
        weight_mem[16'h2B95] <= 0;
        weight_mem[16'h2B96] <= 0;
        weight_mem[16'h2B97] <= 0;
        weight_mem[16'h2B98] <= 0;
        weight_mem[16'h2B99] <= 0;
        weight_mem[16'h2B9A] <= 0;
        weight_mem[16'h2B9B] <= 0;
        weight_mem[16'h2B9C] <= 0;
        weight_mem[16'h2B9D] <= 0;
        weight_mem[16'h2B9E] <= 0;
        weight_mem[16'h2B9F] <= 0;
        weight_mem[16'h2BA0] <= 0;
        weight_mem[16'h2BA1] <= 0;
        weight_mem[16'h2BA2] <= 0;
        weight_mem[16'h2BA3] <= 0;
        weight_mem[16'h2BA4] <= 0;
        weight_mem[16'h2BA5] <= 0;
        weight_mem[16'h2BA6] <= 0;
        weight_mem[16'h2BA7] <= 0;
        weight_mem[16'h2BA8] <= 0;
        weight_mem[16'h2BA9] <= 0;
        weight_mem[16'h2BAA] <= 0;
        weight_mem[16'h2BAB] <= 0;
        weight_mem[16'h2BAC] <= 0;
        weight_mem[16'h2BAD] <= 0;
        weight_mem[16'h2BAE] <= 0;
        weight_mem[16'h2BAF] <= 0;

        // layer 1 neuron 22
        weight_mem[16'h2C00] <= 0;
        weight_mem[16'h2C01] <= 0;
        weight_mem[16'h2C02] <= 0;
        weight_mem[16'h2C03] <= 0;
        weight_mem[16'h2C04] <= 0;
        weight_mem[16'h2C05] <= 0;
        weight_mem[16'h2C06] <= 0;
        weight_mem[16'h2C07] <= 0;
        weight_mem[16'h2C08] <= 0;
        weight_mem[16'h2C09] <= 0;
        weight_mem[16'h2C0A] <= 0;
        weight_mem[16'h2C0B] <= 0;
        weight_mem[16'h2C0C] <= 0;
        weight_mem[16'h2C0D] <= 0;
        weight_mem[16'h2C0E] <= 0;
        weight_mem[16'h2C0F] <= 0;
        weight_mem[16'h2C10] <= 0;
        weight_mem[16'h2C11] <= 0;
        weight_mem[16'h2C12] <= 0;
        weight_mem[16'h2C13] <= 0;
        weight_mem[16'h2C14] <= 0;
        weight_mem[16'h2C15] <= 0;
        weight_mem[16'h2C16] <= 0;
        weight_mem[16'h2C17] <= 0;
        weight_mem[16'h2C18] <= 0;
        weight_mem[16'h2C19] <= 0;
        weight_mem[16'h2C1A] <= 0;
        weight_mem[16'h2C1B] <= 0;
        weight_mem[16'h2C1C] <= 0;
        weight_mem[16'h2C1D] <= 0;
        weight_mem[16'h2C1E] <= 0;
        weight_mem[16'h2C1F] <= 0;
        weight_mem[16'h2C20] <= 0;
        weight_mem[16'h2C21] <= 0;
        weight_mem[16'h2C22] <= 0;
        weight_mem[16'h2C23] <= 0;
        weight_mem[16'h2C24] <= 0;
        weight_mem[16'h2C25] <= 0;
        weight_mem[16'h2C26] <= 0;
        weight_mem[16'h2C27] <= 0;
        weight_mem[16'h2C28] <= 0;
        weight_mem[16'h2C29] <= 0;
        weight_mem[16'h2C2A] <= 0;
        weight_mem[16'h2C2B] <= 0;
        weight_mem[16'h2C2C] <= 0;
        weight_mem[16'h2C2D] <= 0;
        weight_mem[16'h2C2E] <= 0;
        weight_mem[16'h2C2F] <= 0;
        weight_mem[16'h2C30] <= 0;
        weight_mem[16'h2C31] <= 0;
        weight_mem[16'h2C32] <= 0;
        weight_mem[16'h2C33] <= 0;
        weight_mem[16'h2C34] <= 0;
        weight_mem[16'h2C35] <= 0;
        weight_mem[16'h2C36] <= 0;
        weight_mem[16'h2C37] <= 0;
        weight_mem[16'h2C38] <= 0;
        weight_mem[16'h2C39] <= 0;
        weight_mem[16'h2C3A] <= 0;
        weight_mem[16'h2C3B] <= 0;
        weight_mem[16'h2C3C] <= 0;
        weight_mem[16'h2C3D] <= 0;
        weight_mem[16'h2C3E] <= 0;
        weight_mem[16'h2C3F] <= 0;
        weight_mem[16'h2C40] <= 0;
        weight_mem[16'h2C41] <= 0;
        weight_mem[16'h2C42] <= 0;
        weight_mem[16'h2C43] <= 0;
        weight_mem[16'h2C44] <= 0;
        weight_mem[16'h2C45] <= 0;
        weight_mem[16'h2C46] <= 0;
        weight_mem[16'h2C47] <= 0;
        weight_mem[16'h2C48] <= 0;
        weight_mem[16'h2C49] <= 0;
        weight_mem[16'h2C4A] <= 0;
        weight_mem[16'h2C4B] <= 0;
        weight_mem[16'h2C4C] <= 0;
        weight_mem[16'h2C4D] <= 0;
        weight_mem[16'h2C4E] <= 0;
        weight_mem[16'h2C4F] <= 0;
        weight_mem[16'h2C50] <= 0;
        weight_mem[16'h2C51] <= 0;
        weight_mem[16'h2C52] <= 0;
        weight_mem[16'h2C53] <= 0;
        weight_mem[16'h2C54] <= 0;
        weight_mem[16'h2C55] <= 0;
        weight_mem[16'h2C56] <= 0;
        weight_mem[16'h2C57] <= 0;
        weight_mem[16'h2C58] <= 0;
        weight_mem[16'h2C59] <= 0;
        weight_mem[16'h2C5A] <= 0;
        weight_mem[16'h2C5B] <= 0;
        weight_mem[16'h2C5C] <= 0;
        weight_mem[16'h2C5D] <= 0;
        weight_mem[16'h2C5E] <= 0;
        weight_mem[16'h2C5F] <= 0;
        weight_mem[16'h2C60] <= 0;
        weight_mem[16'h2C61] <= 0;
        weight_mem[16'h2C62] <= 0;
        weight_mem[16'h2C63] <= 0;
        weight_mem[16'h2C64] <= 0;
        weight_mem[16'h2C65] <= 0;
        weight_mem[16'h2C66] <= 0;
        weight_mem[16'h2C67] <= 0;
        weight_mem[16'h2C68] <= 0;
        weight_mem[16'h2C69] <= 0;
        weight_mem[16'h2C6A] <= 0;
        weight_mem[16'h2C6B] <= 0;
        weight_mem[16'h2C6C] <= 0;
        weight_mem[16'h2C6D] <= 0;
        weight_mem[16'h2C6E] <= 0;
        weight_mem[16'h2C6F] <= 0;
        weight_mem[16'h2C70] <= 0;
        weight_mem[16'h2C71] <= 0;
        weight_mem[16'h2C72] <= 0;
        weight_mem[16'h2C73] <= 0;
        weight_mem[16'h2C74] <= 0;
        weight_mem[16'h2C75] <= 0;
        weight_mem[16'h2C76] <= 0;
        weight_mem[16'h2C77] <= 0;
        weight_mem[16'h2C78] <= 0;
        weight_mem[16'h2C79] <= 0;
        weight_mem[16'h2C7A] <= 0;
        weight_mem[16'h2C7B] <= 0;
        weight_mem[16'h2C7C] <= 0;
        weight_mem[16'h2C7D] <= 0;
        weight_mem[16'h2C7E] <= 0;
        weight_mem[16'h2C7F] <= 0;
        weight_mem[16'h2C80] <= 0;
        weight_mem[16'h2C81] <= 0;
        weight_mem[16'h2C82] <= 0;
        weight_mem[16'h2C83] <= 0;
        weight_mem[16'h2C84] <= 0;
        weight_mem[16'h2C85] <= 0;
        weight_mem[16'h2C86] <= 0;
        weight_mem[16'h2C87] <= 0;
        weight_mem[16'h2C88] <= 0;
        weight_mem[16'h2C89] <= 0;
        weight_mem[16'h2C8A] <= 0;
        weight_mem[16'h2C8B] <= 0;
        weight_mem[16'h2C8C] <= 0;
        weight_mem[16'h2C8D] <= 0;
        weight_mem[16'h2C8E] <= 0;
        weight_mem[16'h2C8F] <= 0;
        weight_mem[16'h2C90] <= 0;
        weight_mem[16'h2C91] <= 0;
        weight_mem[16'h2C92] <= 0;
        weight_mem[16'h2C93] <= 0;
        weight_mem[16'h2C94] <= 0;
        weight_mem[16'h2C95] <= 0;
        weight_mem[16'h2C96] <= 0;
        weight_mem[16'h2C97] <= 0;
        weight_mem[16'h2C98] <= 0;
        weight_mem[16'h2C99] <= 0;
        weight_mem[16'h2C9A] <= 0;
        weight_mem[16'h2C9B] <= 0;
        weight_mem[16'h2C9C] <= 0;
        weight_mem[16'h2C9D] <= 0;
        weight_mem[16'h2C9E] <= 0;
        weight_mem[16'h2C9F] <= 0;
        weight_mem[16'h2CA0] <= 0;
        weight_mem[16'h2CA1] <= 0;
        weight_mem[16'h2CA2] <= 0;
        weight_mem[16'h2CA3] <= 0;
        weight_mem[16'h2CA4] <= 0;
        weight_mem[16'h2CA5] <= 0;
        weight_mem[16'h2CA6] <= 0;
        weight_mem[16'h2CA7] <= 0;
        weight_mem[16'h2CA8] <= 0;
        weight_mem[16'h2CA9] <= 0;
        weight_mem[16'h2CAA] <= 0;
        weight_mem[16'h2CAB] <= 0;
        weight_mem[16'h2CAC] <= 0;
        weight_mem[16'h2CAD] <= 0;
        weight_mem[16'h2CAE] <= 0;
        weight_mem[16'h2CAF] <= 0;
        weight_mem[16'h2CB0] <= 0;
        weight_mem[16'h2CB1] <= 0;
        weight_mem[16'h2CB2] <= 0;
        weight_mem[16'h2CB3] <= 0;
        weight_mem[16'h2CB4] <= 0;
        weight_mem[16'h2CB5] <= 0;
        weight_mem[16'h2CB6] <= 0;
        weight_mem[16'h2CB7] <= 0;
        weight_mem[16'h2CB8] <= 0;
        weight_mem[16'h2CB9] <= 0;
        weight_mem[16'h2CBA] <= 0;
        weight_mem[16'h2CBB] <= 0;
        weight_mem[16'h2CBC] <= 0;
        weight_mem[16'h2CBD] <= 0;
        weight_mem[16'h2CBE] <= 0;
        weight_mem[16'h2CBF] <= 0;
        weight_mem[16'h2CC0] <= 0;
        weight_mem[16'h2CC1] <= 0;
        weight_mem[16'h2CC2] <= 0;
        weight_mem[16'h2CC3] <= 0;
        weight_mem[16'h2CC4] <= 0;
        weight_mem[16'h2CC5] <= 0;
        weight_mem[16'h2CC6] <= 0;
        weight_mem[16'h2CC7] <= 0;
        weight_mem[16'h2CC8] <= 0;
        weight_mem[16'h2CC9] <= 0;
        weight_mem[16'h2CCA] <= 0;
        weight_mem[16'h2CCB] <= 0;
        weight_mem[16'h2CCC] <= 0;
        weight_mem[16'h2CCD] <= 0;
        weight_mem[16'h2CCE] <= 0;
        weight_mem[16'h2CCF] <= 0;
        weight_mem[16'h2CD0] <= 0;
        weight_mem[16'h2CD1] <= 0;
        weight_mem[16'h2CD2] <= 0;
        weight_mem[16'h2CD3] <= 0;
        weight_mem[16'h2CD4] <= 0;
        weight_mem[16'h2CD5] <= 0;
        weight_mem[16'h2CD6] <= 0;
        weight_mem[16'h2CD7] <= 0;
        weight_mem[16'h2CD8] <= 0;
        weight_mem[16'h2CD9] <= 0;
        weight_mem[16'h2CDA] <= 0;
        weight_mem[16'h2CDB] <= 0;
        weight_mem[16'h2CDC] <= 0;
        weight_mem[16'h2CDD] <= 0;
        weight_mem[16'h2CDE] <= 0;
        weight_mem[16'h2CDF] <= 0;
        weight_mem[16'h2CE0] <= 0;
        weight_mem[16'h2CE1] <= 0;
        weight_mem[16'h2CE2] <= 0;
        weight_mem[16'h2CE3] <= 0;
        weight_mem[16'h2CE4] <= 0;
        weight_mem[16'h2CE5] <= 0;
        weight_mem[16'h2CE6] <= 0;
        weight_mem[16'h2CE7] <= 0;
        weight_mem[16'h2CE8] <= 0;
        weight_mem[16'h2CE9] <= 0;
        weight_mem[16'h2CEA] <= 0;
        weight_mem[16'h2CEB] <= 0;
        weight_mem[16'h2CEC] <= 0;
        weight_mem[16'h2CED] <= 0;
        weight_mem[16'h2CEE] <= 0;
        weight_mem[16'h2CEF] <= 0;
        weight_mem[16'h2CF0] <= 0;
        weight_mem[16'h2CF1] <= 0;
        weight_mem[16'h2CF2] <= 0;
        weight_mem[16'h2CF3] <= 0;
        weight_mem[16'h2CF4] <= 0;
        weight_mem[16'h2CF5] <= 0;
        weight_mem[16'h2CF6] <= 0;
        weight_mem[16'h2CF7] <= 0;
        weight_mem[16'h2CF8] <= 0;
        weight_mem[16'h2CF9] <= 0;
        weight_mem[16'h2CFA] <= 0;
        weight_mem[16'h2CFB] <= 0;
        weight_mem[16'h2CFC] <= 0;
        weight_mem[16'h2CFD] <= 0;
        weight_mem[16'h2CFE] <= 0;
        weight_mem[16'h2CFF] <= 0;
        weight_mem[16'h2D00] <= 0;
        weight_mem[16'h2D01] <= 0;
        weight_mem[16'h2D02] <= 0;
        weight_mem[16'h2D03] <= 0;
        weight_mem[16'h2D04] <= 0;
        weight_mem[16'h2D05] <= 0;
        weight_mem[16'h2D06] <= 0;
        weight_mem[16'h2D07] <= 0;
        weight_mem[16'h2D08] <= 0;
        weight_mem[16'h2D09] <= 0;
        weight_mem[16'h2D0A] <= 0;
        weight_mem[16'h2D0B] <= 0;
        weight_mem[16'h2D0C] <= 0;
        weight_mem[16'h2D0D] <= 0;
        weight_mem[16'h2D0E] <= 0;
        weight_mem[16'h2D0F] <= 0;
        weight_mem[16'h2D10] <= 0;
        weight_mem[16'h2D11] <= 0;
        weight_mem[16'h2D12] <= 0;
        weight_mem[16'h2D13] <= 0;
        weight_mem[16'h2D14] <= 0;
        weight_mem[16'h2D15] <= 0;
        weight_mem[16'h2D16] <= 0;
        weight_mem[16'h2D17] <= 0;
        weight_mem[16'h2D18] <= 0;
        weight_mem[16'h2D19] <= 0;
        weight_mem[16'h2D1A] <= 0;
        weight_mem[16'h2D1B] <= 0;
        weight_mem[16'h2D1C] <= 0;
        weight_mem[16'h2D1D] <= 0;
        weight_mem[16'h2D1E] <= 0;
        weight_mem[16'h2D1F] <= 0;
        weight_mem[16'h2D20] <= 0;
        weight_mem[16'h2D21] <= 0;
        weight_mem[16'h2D22] <= 0;
        weight_mem[16'h2D23] <= 0;
        weight_mem[16'h2D24] <= 0;
        weight_mem[16'h2D25] <= 0;
        weight_mem[16'h2D26] <= 0;
        weight_mem[16'h2D27] <= 0;
        weight_mem[16'h2D28] <= 0;
        weight_mem[16'h2D29] <= 0;
        weight_mem[16'h2D2A] <= 0;
        weight_mem[16'h2D2B] <= 0;
        weight_mem[16'h2D2C] <= 0;
        weight_mem[16'h2D2D] <= 0;
        weight_mem[16'h2D2E] <= 0;
        weight_mem[16'h2D2F] <= 0;
        weight_mem[16'h2D30] <= 0;
        weight_mem[16'h2D31] <= 0;
        weight_mem[16'h2D32] <= 0;
        weight_mem[16'h2D33] <= 0;
        weight_mem[16'h2D34] <= 0;
        weight_mem[16'h2D35] <= 0;
        weight_mem[16'h2D36] <= 0;
        weight_mem[16'h2D37] <= 0;
        weight_mem[16'h2D38] <= 0;
        weight_mem[16'h2D39] <= 0;
        weight_mem[16'h2D3A] <= 0;
        weight_mem[16'h2D3B] <= 0;
        weight_mem[16'h2D3C] <= 0;
        weight_mem[16'h2D3D] <= 0;
        weight_mem[16'h2D3E] <= 0;
        weight_mem[16'h2D3F] <= 0;
        weight_mem[16'h2D40] <= 0;
        weight_mem[16'h2D41] <= 0;
        weight_mem[16'h2D42] <= 0;
        weight_mem[16'h2D43] <= 0;
        weight_mem[16'h2D44] <= 0;
        weight_mem[16'h2D45] <= 0;
        weight_mem[16'h2D46] <= 0;
        weight_mem[16'h2D47] <= 0;
        weight_mem[16'h2D48] <= 0;
        weight_mem[16'h2D49] <= 0;
        weight_mem[16'h2D4A] <= 0;
        weight_mem[16'h2D4B] <= 0;
        weight_mem[16'h2D4C] <= 0;
        weight_mem[16'h2D4D] <= 0;
        weight_mem[16'h2D4E] <= 0;
        weight_mem[16'h2D4F] <= 0;
        weight_mem[16'h2D50] <= 0;
        weight_mem[16'h2D51] <= 0;
        weight_mem[16'h2D52] <= 0;
        weight_mem[16'h2D53] <= 0;
        weight_mem[16'h2D54] <= 0;
        weight_mem[16'h2D55] <= 0;
        weight_mem[16'h2D56] <= 0;
        weight_mem[16'h2D57] <= 0;
        weight_mem[16'h2D58] <= 0;
        weight_mem[16'h2D59] <= 0;
        weight_mem[16'h2D5A] <= 0;
        weight_mem[16'h2D5B] <= 0;
        weight_mem[16'h2D5C] <= 0;
        weight_mem[16'h2D5D] <= 0;
        weight_mem[16'h2D5E] <= 0;
        weight_mem[16'h2D5F] <= 0;
        weight_mem[16'h2D60] <= 0;
        weight_mem[16'h2D61] <= 0;
        weight_mem[16'h2D62] <= 0;
        weight_mem[16'h2D63] <= 0;
        weight_mem[16'h2D64] <= 0;
        weight_mem[16'h2D65] <= 0;
        weight_mem[16'h2D66] <= 0;
        weight_mem[16'h2D67] <= 0;
        weight_mem[16'h2D68] <= 0;
        weight_mem[16'h2D69] <= 0;
        weight_mem[16'h2D6A] <= 0;
        weight_mem[16'h2D6B] <= 0;
        weight_mem[16'h2D6C] <= 0;
        weight_mem[16'h2D6D] <= 0;
        weight_mem[16'h2D6E] <= 0;
        weight_mem[16'h2D6F] <= 0;
        weight_mem[16'h2D70] <= 0;
        weight_mem[16'h2D71] <= 0;
        weight_mem[16'h2D72] <= 0;
        weight_mem[16'h2D73] <= 0;
        weight_mem[16'h2D74] <= 0;
        weight_mem[16'h2D75] <= 0;
        weight_mem[16'h2D76] <= 0;
        weight_mem[16'h2D77] <= 0;
        weight_mem[16'h2D78] <= 0;
        weight_mem[16'h2D79] <= 0;
        weight_mem[16'h2D7A] <= 0;
        weight_mem[16'h2D7B] <= 0;
        weight_mem[16'h2D7C] <= 0;
        weight_mem[16'h2D7D] <= 0;
        weight_mem[16'h2D7E] <= 0;
        weight_mem[16'h2D7F] <= 0;
        weight_mem[16'h2D80] <= 0;
        weight_mem[16'h2D81] <= 0;
        weight_mem[16'h2D82] <= 0;
        weight_mem[16'h2D83] <= 0;
        weight_mem[16'h2D84] <= 0;
        weight_mem[16'h2D85] <= 0;
        weight_mem[16'h2D86] <= 0;
        weight_mem[16'h2D87] <= 0;
        weight_mem[16'h2D88] <= 0;
        weight_mem[16'h2D89] <= 0;
        weight_mem[16'h2D8A] <= 0;
        weight_mem[16'h2D8B] <= 0;
        weight_mem[16'h2D8C] <= 0;
        weight_mem[16'h2D8D] <= 0;
        weight_mem[16'h2D8E] <= 0;
        weight_mem[16'h2D8F] <= 0;
        weight_mem[16'h2D90] <= 0;
        weight_mem[16'h2D91] <= 0;
        weight_mem[16'h2D92] <= 0;
        weight_mem[16'h2D93] <= 0;
        weight_mem[16'h2D94] <= 0;
        weight_mem[16'h2D95] <= 0;
        weight_mem[16'h2D96] <= 0;
        weight_mem[16'h2D97] <= 0;
        weight_mem[16'h2D98] <= 0;
        weight_mem[16'h2D99] <= 0;
        weight_mem[16'h2D9A] <= 0;
        weight_mem[16'h2D9B] <= 0;
        weight_mem[16'h2D9C] <= 0;
        weight_mem[16'h2D9D] <= 0;
        weight_mem[16'h2D9E] <= 0;
        weight_mem[16'h2D9F] <= 0;
        weight_mem[16'h2DA0] <= 0;
        weight_mem[16'h2DA1] <= 0;
        weight_mem[16'h2DA2] <= 0;
        weight_mem[16'h2DA3] <= 0;
        weight_mem[16'h2DA4] <= 0;
        weight_mem[16'h2DA5] <= 0;
        weight_mem[16'h2DA6] <= 0;
        weight_mem[16'h2DA7] <= 0;
        weight_mem[16'h2DA8] <= 0;
        weight_mem[16'h2DA9] <= 0;
        weight_mem[16'h2DAA] <= 0;
        weight_mem[16'h2DAB] <= 0;
        weight_mem[16'h2DAC] <= 0;
        weight_mem[16'h2DAD] <= 0;
        weight_mem[16'h2DAE] <= 0;
        weight_mem[16'h2DAF] <= 0;

        // layer 1 neuron 23
        weight_mem[16'h2E00] <= 0;
        weight_mem[16'h2E01] <= 0;
        weight_mem[16'h2E02] <= 0;
        weight_mem[16'h2E03] <= 0;
        weight_mem[16'h2E04] <= 0;
        weight_mem[16'h2E05] <= 0;
        weight_mem[16'h2E06] <= 0;
        weight_mem[16'h2E07] <= 0;
        weight_mem[16'h2E08] <= 0;
        weight_mem[16'h2E09] <= 0;
        weight_mem[16'h2E0A] <= 0;
        weight_mem[16'h2E0B] <= 0;
        weight_mem[16'h2E0C] <= 0;
        weight_mem[16'h2E0D] <= 0;
        weight_mem[16'h2E0E] <= 0;
        weight_mem[16'h2E0F] <= 0;
        weight_mem[16'h2E10] <= 0;
        weight_mem[16'h2E11] <= 0;
        weight_mem[16'h2E12] <= 0;
        weight_mem[16'h2E13] <= 0;
        weight_mem[16'h2E14] <= 0;
        weight_mem[16'h2E15] <= 0;
        weight_mem[16'h2E16] <= 0;
        weight_mem[16'h2E17] <= 0;
        weight_mem[16'h2E18] <= 0;
        weight_mem[16'h2E19] <= 0;
        weight_mem[16'h2E1A] <= 0;
        weight_mem[16'h2E1B] <= 0;
        weight_mem[16'h2E1C] <= 0;
        weight_mem[16'h2E1D] <= 0;
        weight_mem[16'h2E1E] <= 0;
        weight_mem[16'h2E1F] <= 0;
        weight_mem[16'h2E20] <= 0;
        weight_mem[16'h2E21] <= 0;
        weight_mem[16'h2E22] <= 0;
        weight_mem[16'h2E23] <= 0;
        weight_mem[16'h2E24] <= 0;
        weight_mem[16'h2E25] <= 0;
        weight_mem[16'h2E26] <= 0;
        weight_mem[16'h2E27] <= 0;
        weight_mem[16'h2E28] <= 0;
        weight_mem[16'h2E29] <= 0;
        weight_mem[16'h2E2A] <= 0;
        weight_mem[16'h2E2B] <= 0;
        weight_mem[16'h2E2C] <= 0;
        weight_mem[16'h2E2D] <= 0;
        weight_mem[16'h2E2E] <= 0;
        weight_mem[16'h2E2F] <= 0;
        weight_mem[16'h2E30] <= 0;
        weight_mem[16'h2E31] <= 0;
        weight_mem[16'h2E32] <= 0;
        weight_mem[16'h2E33] <= 0;
        weight_mem[16'h2E34] <= 0;
        weight_mem[16'h2E35] <= 0;
        weight_mem[16'h2E36] <= 0;
        weight_mem[16'h2E37] <= 0;
        weight_mem[16'h2E38] <= 0;
        weight_mem[16'h2E39] <= 0;
        weight_mem[16'h2E3A] <= 0;
        weight_mem[16'h2E3B] <= 0;
        weight_mem[16'h2E3C] <= 0;
        weight_mem[16'h2E3D] <= 0;
        weight_mem[16'h2E3E] <= 0;
        weight_mem[16'h2E3F] <= 0;
        weight_mem[16'h2E40] <= 0;
        weight_mem[16'h2E41] <= 0;
        weight_mem[16'h2E42] <= 0;
        weight_mem[16'h2E43] <= 0;
        weight_mem[16'h2E44] <= 0;
        weight_mem[16'h2E45] <= 0;
        weight_mem[16'h2E46] <= 0;
        weight_mem[16'h2E47] <= 0;
        weight_mem[16'h2E48] <= 0;
        weight_mem[16'h2E49] <= 0;
        weight_mem[16'h2E4A] <= 0;
        weight_mem[16'h2E4B] <= 0;
        weight_mem[16'h2E4C] <= 0;
        weight_mem[16'h2E4D] <= 0;
        weight_mem[16'h2E4E] <= 0;
        weight_mem[16'h2E4F] <= 0;
        weight_mem[16'h2E50] <= 0;
        weight_mem[16'h2E51] <= 0;
        weight_mem[16'h2E52] <= 0;
        weight_mem[16'h2E53] <= 0;
        weight_mem[16'h2E54] <= 0;
        weight_mem[16'h2E55] <= 0;
        weight_mem[16'h2E56] <= 0;
        weight_mem[16'h2E57] <= 0;
        weight_mem[16'h2E58] <= 0;
        weight_mem[16'h2E59] <= 0;
        weight_mem[16'h2E5A] <= 0;
        weight_mem[16'h2E5B] <= 0;
        weight_mem[16'h2E5C] <= 0;
        weight_mem[16'h2E5D] <= 0;
        weight_mem[16'h2E5E] <= 0;
        weight_mem[16'h2E5F] <= 0;
        weight_mem[16'h2E60] <= 0;
        weight_mem[16'h2E61] <= 0;
        weight_mem[16'h2E62] <= 0;
        weight_mem[16'h2E63] <= 0;
        weight_mem[16'h2E64] <= 0;
        weight_mem[16'h2E65] <= 0;
        weight_mem[16'h2E66] <= 0;
        weight_mem[16'h2E67] <= 0;
        weight_mem[16'h2E68] <= 0;
        weight_mem[16'h2E69] <= 0;
        weight_mem[16'h2E6A] <= 0;
        weight_mem[16'h2E6B] <= 0;
        weight_mem[16'h2E6C] <= 0;
        weight_mem[16'h2E6D] <= 0;
        weight_mem[16'h2E6E] <= 0;
        weight_mem[16'h2E6F] <= 0;
        weight_mem[16'h2E70] <= 0;
        weight_mem[16'h2E71] <= 0;
        weight_mem[16'h2E72] <= 0;
        weight_mem[16'h2E73] <= 0;
        weight_mem[16'h2E74] <= 0;
        weight_mem[16'h2E75] <= 0;
        weight_mem[16'h2E76] <= 0;
        weight_mem[16'h2E77] <= 0;
        weight_mem[16'h2E78] <= 0;
        weight_mem[16'h2E79] <= 0;
        weight_mem[16'h2E7A] <= 0;
        weight_mem[16'h2E7B] <= 0;
        weight_mem[16'h2E7C] <= 0;
        weight_mem[16'h2E7D] <= 0;
        weight_mem[16'h2E7E] <= 0;
        weight_mem[16'h2E7F] <= 0;
        weight_mem[16'h2E80] <= 0;
        weight_mem[16'h2E81] <= 0;
        weight_mem[16'h2E82] <= 0;
        weight_mem[16'h2E83] <= 0;
        weight_mem[16'h2E84] <= 0;
        weight_mem[16'h2E85] <= 0;
        weight_mem[16'h2E86] <= 0;
        weight_mem[16'h2E87] <= 0;
        weight_mem[16'h2E88] <= 0;
        weight_mem[16'h2E89] <= 0;
        weight_mem[16'h2E8A] <= 0;
        weight_mem[16'h2E8B] <= 0;
        weight_mem[16'h2E8C] <= 0;
        weight_mem[16'h2E8D] <= 0;
        weight_mem[16'h2E8E] <= 0;
        weight_mem[16'h2E8F] <= 0;
        weight_mem[16'h2E90] <= 0;
        weight_mem[16'h2E91] <= 0;
        weight_mem[16'h2E92] <= 0;
        weight_mem[16'h2E93] <= 0;
        weight_mem[16'h2E94] <= 0;
        weight_mem[16'h2E95] <= 0;
        weight_mem[16'h2E96] <= 0;
        weight_mem[16'h2E97] <= 0;
        weight_mem[16'h2E98] <= 0;
        weight_mem[16'h2E99] <= 0;
        weight_mem[16'h2E9A] <= 0;
        weight_mem[16'h2E9B] <= 0;
        weight_mem[16'h2E9C] <= 0;
        weight_mem[16'h2E9D] <= 0;
        weight_mem[16'h2E9E] <= 0;
        weight_mem[16'h2E9F] <= 0;
        weight_mem[16'h2EA0] <= 0;
        weight_mem[16'h2EA1] <= 0;
        weight_mem[16'h2EA2] <= 0;
        weight_mem[16'h2EA3] <= 0;
        weight_mem[16'h2EA4] <= 0;
        weight_mem[16'h2EA5] <= 0;
        weight_mem[16'h2EA6] <= 0;
        weight_mem[16'h2EA7] <= 0;
        weight_mem[16'h2EA8] <= 0;
        weight_mem[16'h2EA9] <= 0;
        weight_mem[16'h2EAA] <= 0;
        weight_mem[16'h2EAB] <= 0;
        weight_mem[16'h2EAC] <= 0;
        weight_mem[16'h2EAD] <= 0;
        weight_mem[16'h2EAE] <= 0;
        weight_mem[16'h2EAF] <= 0;
        weight_mem[16'h2EB0] <= 0;
        weight_mem[16'h2EB1] <= 0;
        weight_mem[16'h2EB2] <= 0;
        weight_mem[16'h2EB3] <= 0;
        weight_mem[16'h2EB4] <= 0;
        weight_mem[16'h2EB5] <= 0;
        weight_mem[16'h2EB6] <= 0;
        weight_mem[16'h2EB7] <= 0;
        weight_mem[16'h2EB8] <= 0;
        weight_mem[16'h2EB9] <= 0;
        weight_mem[16'h2EBA] <= 0;
        weight_mem[16'h2EBB] <= 0;
        weight_mem[16'h2EBC] <= 0;
        weight_mem[16'h2EBD] <= 0;
        weight_mem[16'h2EBE] <= 0;
        weight_mem[16'h2EBF] <= 0;
        weight_mem[16'h2EC0] <= 0;
        weight_mem[16'h2EC1] <= 0;
        weight_mem[16'h2EC2] <= 0;
        weight_mem[16'h2EC3] <= 0;
        weight_mem[16'h2EC4] <= 0;
        weight_mem[16'h2EC5] <= 0;
        weight_mem[16'h2EC6] <= 0;
        weight_mem[16'h2EC7] <= 0;
        weight_mem[16'h2EC8] <= 0;
        weight_mem[16'h2EC9] <= 0;
        weight_mem[16'h2ECA] <= 0;
        weight_mem[16'h2ECB] <= 0;
        weight_mem[16'h2ECC] <= 0;
        weight_mem[16'h2ECD] <= 0;
        weight_mem[16'h2ECE] <= 0;
        weight_mem[16'h2ECF] <= 0;
        weight_mem[16'h2ED0] <= 0;
        weight_mem[16'h2ED1] <= 0;
        weight_mem[16'h2ED2] <= 0;
        weight_mem[16'h2ED3] <= 0;
        weight_mem[16'h2ED4] <= 0;
        weight_mem[16'h2ED5] <= 0;
        weight_mem[16'h2ED6] <= 0;
        weight_mem[16'h2ED7] <= 0;
        weight_mem[16'h2ED8] <= 0;
        weight_mem[16'h2ED9] <= 0;
        weight_mem[16'h2EDA] <= 0;
        weight_mem[16'h2EDB] <= 0;
        weight_mem[16'h2EDC] <= 0;
        weight_mem[16'h2EDD] <= 0;
        weight_mem[16'h2EDE] <= 0;
        weight_mem[16'h2EDF] <= 0;
        weight_mem[16'h2EE0] <= 0;
        weight_mem[16'h2EE1] <= 0;
        weight_mem[16'h2EE2] <= 0;
        weight_mem[16'h2EE3] <= 0;
        weight_mem[16'h2EE4] <= 0;
        weight_mem[16'h2EE5] <= 0;
        weight_mem[16'h2EE6] <= 0;
        weight_mem[16'h2EE7] <= 0;
        weight_mem[16'h2EE8] <= 0;
        weight_mem[16'h2EE9] <= 0;
        weight_mem[16'h2EEA] <= 0;
        weight_mem[16'h2EEB] <= 0;
        weight_mem[16'h2EEC] <= 0;
        weight_mem[16'h2EED] <= 0;
        weight_mem[16'h2EEE] <= 0;
        weight_mem[16'h2EEF] <= 0;
        weight_mem[16'h2EF0] <= 0;
        weight_mem[16'h2EF1] <= 0;
        weight_mem[16'h2EF2] <= 0;
        weight_mem[16'h2EF3] <= 0;
        weight_mem[16'h2EF4] <= 0;
        weight_mem[16'h2EF5] <= 0;
        weight_mem[16'h2EF6] <= 0;
        weight_mem[16'h2EF7] <= 0;
        weight_mem[16'h2EF8] <= 0;
        weight_mem[16'h2EF9] <= 0;
        weight_mem[16'h2EFA] <= 0;
        weight_mem[16'h2EFB] <= 0;
        weight_mem[16'h2EFC] <= 0;
        weight_mem[16'h2EFD] <= 0;
        weight_mem[16'h2EFE] <= 0;
        weight_mem[16'h2EFF] <= 0;
        weight_mem[16'h2F00] <= 0;
        weight_mem[16'h2F01] <= 0;
        weight_mem[16'h2F02] <= 0;
        weight_mem[16'h2F03] <= 0;
        weight_mem[16'h2F04] <= 0;
        weight_mem[16'h2F05] <= 0;
        weight_mem[16'h2F06] <= 0;
        weight_mem[16'h2F07] <= 0;
        weight_mem[16'h2F08] <= 0;
        weight_mem[16'h2F09] <= 0;
        weight_mem[16'h2F0A] <= 0;
        weight_mem[16'h2F0B] <= 0;
        weight_mem[16'h2F0C] <= 0;
        weight_mem[16'h2F0D] <= 0;
        weight_mem[16'h2F0E] <= 0;
        weight_mem[16'h2F0F] <= 0;
        weight_mem[16'h2F10] <= 0;
        weight_mem[16'h2F11] <= 0;
        weight_mem[16'h2F12] <= 0;
        weight_mem[16'h2F13] <= 0;
        weight_mem[16'h2F14] <= 0;
        weight_mem[16'h2F15] <= 0;
        weight_mem[16'h2F16] <= 0;
        weight_mem[16'h2F17] <= 0;
        weight_mem[16'h2F18] <= 0;
        weight_mem[16'h2F19] <= 0;
        weight_mem[16'h2F1A] <= 0;
        weight_mem[16'h2F1B] <= 0;
        weight_mem[16'h2F1C] <= 0;
        weight_mem[16'h2F1D] <= 0;
        weight_mem[16'h2F1E] <= 0;
        weight_mem[16'h2F1F] <= 0;
        weight_mem[16'h2F20] <= 0;
        weight_mem[16'h2F21] <= 0;
        weight_mem[16'h2F22] <= 0;
        weight_mem[16'h2F23] <= 0;
        weight_mem[16'h2F24] <= 0;
        weight_mem[16'h2F25] <= 0;
        weight_mem[16'h2F26] <= 0;
        weight_mem[16'h2F27] <= 0;
        weight_mem[16'h2F28] <= 0;
        weight_mem[16'h2F29] <= 0;
        weight_mem[16'h2F2A] <= 0;
        weight_mem[16'h2F2B] <= 0;
        weight_mem[16'h2F2C] <= 0;
        weight_mem[16'h2F2D] <= 0;
        weight_mem[16'h2F2E] <= 0;
        weight_mem[16'h2F2F] <= 0;
        weight_mem[16'h2F30] <= 0;
        weight_mem[16'h2F31] <= 0;
        weight_mem[16'h2F32] <= 0;
        weight_mem[16'h2F33] <= 0;
        weight_mem[16'h2F34] <= 0;
        weight_mem[16'h2F35] <= 0;
        weight_mem[16'h2F36] <= 0;
        weight_mem[16'h2F37] <= 0;
        weight_mem[16'h2F38] <= 0;
        weight_mem[16'h2F39] <= 0;
        weight_mem[16'h2F3A] <= 0;
        weight_mem[16'h2F3B] <= 0;
        weight_mem[16'h2F3C] <= 0;
        weight_mem[16'h2F3D] <= 0;
        weight_mem[16'h2F3E] <= 0;
        weight_mem[16'h2F3F] <= 0;
        weight_mem[16'h2F40] <= 0;
        weight_mem[16'h2F41] <= 0;
        weight_mem[16'h2F42] <= 0;
        weight_mem[16'h2F43] <= 0;
        weight_mem[16'h2F44] <= 0;
        weight_mem[16'h2F45] <= 0;
        weight_mem[16'h2F46] <= 0;
        weight_mem[16'h2F47] <= 0;
        weight_mem[16'h2F48] <= 0;
        weight_mem[16'h2F49] <= 0;
        weight_mem[16'h2F4A] <= 0;
        weight_mem[16'h2F4B] <= 0;
        weight_mem[16'h2F4C] <= 0;
        weight_mem[16'h2F4D] <= 0;
        weight_mem[16'h2F4E] <= 0;
        weight_mem[16'h2F4F] <= 0;
        weight_mem[16'h2F50] <= 0;
        weight_mem[16'h2F51] <= 0;
        weight_mem[16'h2F52] <= 0;
        weight_mem[16'h2F53] <= 0;
        weight_mem[16'h2F54] <= 0;
        weight_mem[16'h2F55] <= 0;
        weight_mem[16'h2F56] <= 0;
        weight_mem[16'h2F57] <= 0;
        weight_mem[16'h2F58] <= 0;
        weight_mem[16'h2F59] <= 0;
        weight_mem[16'h2F5A] <= 0;
        weight_mem[16'h2F5B] <= 0;
        weight_mem[16'h2F5C] <= 0;
        weight_mem[16'h2F5D] <= 0;
        weight_mem[16'h2F5E] <= 0;
        weight_mem[16'h2F5F] <= 0;
        weight_mem[16'h2F60] <= 0;
        weight_mem[16'h2F61] <= 0;
        weight_mem[16'h2F62] <= 0;
        weight_mem[16'h2F63] <= 0;
        weight_mem[16'h2F64] <= 0;
        weight_mem[16'h2F65] <= 0;
        weight_mem[16'h2F66] <= 0;
        weight_mem[16'h2F67] <= 0;
        weight_mem[16'h2F68] <= 0;
        weight_mem[16'h2F69] <= 0;
        weight_mem[16'h2F6A] <= 0;
        weight_mem[16'h2F6B] <= 0;
        weight_mem[16'h2F6C] <= 0;
        weight_mem[16'h2F6D] <= 0;
        weight_mem[16'h2F6E] <= 0;
        weight_mem[16'h2F6F] <= 0;
        weight_mem[16'h2F70] <= 0;
        weight_mem[16'h2F71] <= 0;
        weight_mem[16'h2F72] <= 0;
        weight_mem[16'h2F73] <= 0;
        weight_mem[16'h2F74] <= 0;
        weight_mem[16'h2F75] <= 0;
        weight_mem[16'h2F76] <= 0;
        weight_mem[16'h2F77] <= 0;
        weight_mem[16'h2F78] <= 0;
        weight_mem[16'h2F79] <= 0;
        weight_mem[16'h2F7A] <= 0;
        weight_mem[16'h2F7B] <= 0;
        weight_mem[16'h2F7C] <= 0;
        weight_mem[16'h2F7D] <= 0;
        weight_mem[16'h2F7E] <= 0;
        weight_mem[16'h2F7F] <= 0;
        weight_mem[16'h2F80] <= 0;
        weight_mem[16'h2F81] <= 0;
        weight_mem[16'h2F82] <= 0;
        weight_mem[16'h2F83] <= 0;
        weight_mem[16'h2F84] <= 0;
        weight_mem[16'h2F85] <= 0;
        weight_mem[16'h2F86] <= 0;
        weight_mem[16'h2F87] <= 0;
        weight_mem[16'h2F88] <= 0;
        weight_mem[16'h2F89] <= 0;
        weight_mem[16'h2F8A] <= 0;
        weight_mem[16'h2F8B] <= 0;
        weight_mem[16'h2F8C] <= 0;
        weight_mem[16'h2F8D] <= 0;
        weight_mem[16'h2F8E] <= 0;
        weight_mem[16'h2F8F] <= 0;
        weight_mem[16'h2F90] <= 0;
        weight_mem[16'h2F91] <= 0;
        weight_mem[16'h2F92] <= 0;
        weight_mem[16'h2F93] <= 0;
        weight_mem[16'h2F94] <= 0;
        weight_mem[16'h2F95] <= 0;
        weight_mem[16'h2F96] <= 0;
        weight_mem[16'h2F97] <= 0;
        weight_mem[16'h2F98] <= 0;
        weight_mem[16'h2F99] <= 0;
        weight_mem[16'h2F9A] <= 0;
        weight_mem[16'h2F9B] <= 0;
        weight_mem[16'h2F9C] <= 0;
        weight_mem[16'h2F9D] <= 0;
        weight_mem[16'h2F9E] <= 0;
        weight_mem[16'h2F9F] <= 0;
        weight_mem[16'h2FA0] <= 0;
        weight_mem[16'h2FA1] <= 0;
        weight_mem[16'h2FA2] <= 0;
        weight_mem[16'h2FA3] <= 0;
        weight_mem[16'h2FA4] <= 0;
        weight_mem[16'h2FA5] <= 0;
        weight_mem[16'h2FA6] <= 0;
        weight_mem[16'h2FA7] <= 0;
        weight_mem[16'h2FA8] <= 0;
        weight_mem[16'h2FA9] <= 0;
        weight_mem[16'h2FAA] <= 0;
        weight_mem[16'h2FAB] <= 0;
        weight_mem[16'h2FAC] <= 0;
        weight_mem[16'h2FAD] <= 0;
        weight_mem[16'h2FAE] <= 0;
        weight_mem[16'h2FAF] <= 0;

        // layer 1 neuron 24
        weight_mem[16'h3000] <= 0;
        weight_mem[16'h3001] <= 0;
        weight_mem[16'h3002] <= 0;
        weight_mem[16'h3003] <= 0;
        weight_mem[16'h3004] <= 0;
        weight_mem[16'h3005] <= 0;
        weight_mem[16'h3006] <= 0;
        weight_mem[16'h3007] <= 0;
        weight_mem[16'h3008] <= 0;
        weight_mem[16'h3009] <= 0;
        weight_mem[16'h300A] <= 0;
        weight_mem[16'h300B] <= 0;
        weight_mem[16'h300C] <= 0;
        weight_mem[16'h300D] <= 0;
        weight_mem[16'h300E] <= 0;
        weight_mem[16'h300F] <= 0;
        weight_mem[16'h3010] <= 0;
        weight_mem[16'h3011] <= 0;
        weight_mem[16'h3012] <= 0;
        weight_mem[16'h3013] <= 0;
        weight_mem[16'h3014] <= 0;
        weight_mem[16'h3015] <= 0;
        weight_mem[16'h3016] <= 0;
        weight_mem[16'h3017] <= 0;
        weight_mem[16'h3018] <= 0;
        weight_mem[16'h3019] <= 0;
        weight_mem[16'h301A] <= 0;
        weight_mem[16'h301B] <= 0;
        weight_mem[16'h301C] <= 0;
        weight_mem[16'h301D] <= 0;
        weight_mem[16'h301E] <= 0;
        weight_mem[16'h301F] <= 0;
        weight_mem[16'h3020] <= 0;
        weight_mem[16'h3021] <= 0;
        weight_mem[16'h3022] <= 0;
        weight_mem[16'h3023] <= 0;
        weight_mem[16'h3024] <= 0;
        weight_mem[16'h3025] <= 0;
        weight_mem[16'h3026] <= 0;
        weight_mem[16'h3027] <= 0;
        weight_mem[16'h3028] <= 0;
        weight_mem[16'h3029] <= 0;
        weight_mem[16'h302A] <= 0;
        weight_mem[16'h302B] <= 0;
        weight_mem[16'h302C] <= 0;
        weight_mem[16'h302D] <= 0;
        weight_mem[16'h302E] <= 0;
        weight_mem[16'h302F] <= 0;
        weight_mem[16'h3030] <= 0;
        weight_mem[16'h3031] <= 0;
        weight_mem[16'h3032] <= 0;
        weight_mem[16'h3033] <= 0;
        weight_mem[16'h3034] <= 0;
        weight_mem[16'h3035] <= 0;
        weight_mem[16'h3036] <= 0;
        weight_mem[16'h3037] <= 0;
        weight_mem[16'h3038] <= 0;
        weight_mem[16'h3039] <= 0;
        weight_mem[16'h303A] <= 0;
        weight_mem[16'h303B] <= 0;
        weight_mem[16'h303C] <= 0;
        weight_mem[16'h303D] <= 0;
        weight_mem[16'h303E] <= 0;
        weight_mem[16'h303F] <= 0;
        weight_mem[16'h3040] <= 0;
        weight_mem[16'h3041] <= 0;
        weight_mem[16'h3042] <= 0;
        weight_mem[16'h3043] <= 0;
        weight_mem[16'h3044] <= 0;
        weight_mem[16'h3045] <= 0;
        weight_mem[16'h3046] <= 0;
        weight_mem[16'h3047] <= 0;
        weight_mem[16'h3048] <= 0;
        weight_mem[16'h3049] <= 0;
        weight_mem[16'h304A] <= 0;
        weight_mem[16'h304B] <= 0;
        weight_mem[16'h304C] <= 0;
        weight_mem[16'h304D] <= 0;
        weight_mem[16'h304E] <= 0;
        weight_mem[16'h304F] <= 0;
        weight_mem[16'h3050] <= 0;
        weight_mem[16'h3051] <= 0;
        weight_mem[16'h3052] <= 0;
        weight_mem[16'h3053] <= 0;
        weight_mem[16'h3054] <= 0;
        weight_mem[16'h3055] <= 0;
        weight_mem[16'h3056] <= 0;
        weight_mem[16'h3057] <= 0;
        weight_mem[16'h3058] <= 0;
        weight_mem[16'h3059] <= 0;
        weight_mem[16'h305A] <= 0;
        weight_mem[16'h305B] <= 0;
        weight_mem[16'h305C] <= 0;
        weight_mem[16'h305D] <= 0;
        weight_mem[16'h305E] <= 0;
        weight_mem[16'h305F] <= 0;
        weight_mem[16'h3060] <= 0;
        weight_mem[16'h3061] <= 0;
        weight_mem[16'h3062] <= 0;
        weight_mem[16'h3063] <= 0;
        weight_mem[16'h3064] <= 0;
        weight_mem[16'h3065] <= 0;
        weight_mem[16'h3066] <= 0;
        weight_mem[16'h3067] <= 0;
        weight_mem[16'h3068] <= 0;
        weight_mem[16'h3069] <= 0;
        weight_mem[16'h306A] <= 0;
        weight_mem[16'h306B] <= 0;
        weight_mem[16'h306C] <= 0;
        weight_mem[16'h306D] <= 0;
        weight_mem[16'h306E] <= 0;
        weight_mem[16'h306F] <= 0;
        weight_mem[16'h3070] <= 0;
        weight_mem[16'h3071] <= 0;
        weight_mem[16'h3072] <= 0;
        weight_mem[16'h3073] <= 0;
        weight_mem[16'h3074] <= 0;
        weight_mem[16'h3075] <= 0;
        weight_mem[16'h3076] <= 0;
        weight_mem[16'h3077] <= 0;
        weight_mem[16'h3078] <= 0;
        weight_mem[16'h3079] <= 0;
        weight_mem[16'h307A] <= 0;
        weight_mem[16'h307B] <= 0;
        weight_mem[16'h307C] <= 0;
        weight_mem[16'h307D] <= 0;
        weight_mem[16'h307E] <= 0;
        weight_mem[16'h307F] <= 0;
        weight_mem[16'h3080] <= 0;
        weight_mem[16'h3081] <= 0;
        weight_mem[16'h3082] <= 0;
        weight_mem[16'h3083] <= 0;
        weight_mem[16'h3084] <= 0;
        weight_mem[16'h3085] <= 0;
        weight_mem[16'h3086] <= 0;
        weight_mem[16'h3087] <= 0;
        weight_mem[16'h3088] <= 0;
        weight_mem[16'h3089] <= 0;
        weight_mem[16'h308A] <= 0;
        weight_mem[16'h308B] <= 0;
        weight_mem[16'h308C] <= 0;
        weight_mem[16'h308D] <= 0;
        weight_mem[16'h308E] <= 0;
        weight_mem[16'h308F] <= 0;
        weight_mem[16'h3090] <= 0;
        weight_mem[16'h3091] <= 0;
        weight_mem[16'h3092] <= 0;
        weight_mem[16'h3093] <= 0;
        weight_mem[16'h3094] <= 0;
        weight_mem[16'h3095] <= 0;
        weight_mem[16'h3096] <= 0;
        weight_mem[16'h3097] <= 0;
        weight_mem[16'h3098] <= 0;
        weight_mem[16'h3099] <= 0;
        weight_mem[16'h309A] <= 0;
        weight_mem[16'h309B] <= 0;
        weight_mem[16'h309C] <= 0;
        weight_mem[16'h309D] <= 0;
        weight_mem[16'h309E] <= 0;
        weight_mem[16'h309F] <= 0;
        weight_mem[16'h30A0] <= 0;
        weight_mem[16'h30A1] <= 0;
        weight_mem[16'h30A2] <= 0;
        weight_mem[16'h30A3] <= 0;
        weight_mem[16'h30A4] <= 0;
        weight_mem[16'h30A5] <= 0;
        weight_mem[16'h30A6] <= 0;
        weight_mem[16'h30A7] <= 0;
        weight_mem[16'h30A8] <= 0;
        weight_mem[16'h30A9] <= 0;
        weight_mem[16'h30AA] <= 0;
        weight_mem[16'h30AB] <= 0;
        weight_mem[16'h30AC] <= 0;
        weight_mem[16'h30AD] <= 0;
        weight_mem[16'h30AE] <= 0;
        weight_mem[16'h30AF] <= 0;
        weight_mem[16'h30B0] <= 0;
        weight_mem[16'h30B1] <= 0;
        weight_mem[16'h30B2] <= 0;
        weight_mem[16'h30B3] <= 0;
        weight_mem[16'h30B4] <= 0;
        weight_mem[16'h30B5] <= 0;
        weight_mem[16'h30B6] <= 0;
        weight_mem[16'h30B7] <= 0;
        weight_mem[16'h30B8] <= 0;
        weight_mem[16'h30B9] <= 0;
        weight_mem[16'h30BA] <= 0;
        weight_mem[16'h30BB] <= 0;
        weight_mem[16'h30BC] <= 0;
        weight_mem[16'h30BD] <= 0;
        weight_mem[16'h30BE] <= 0;
        weight_mem[16'h30BF] <= 0;
        weight_mem[16'h30C0] <= 0;
        weight_mem[16'h30C1] <= 0;
        weight_mem[16'h30C2] <= 0;
        weight_mem[16'h30C3] <= 0;
        weight_mem[16'h30C4] <= 0;
        weight_mem[16'h30C5] <= 0;
        weight_mem[16'h30C6] <= 0;
        weight_mem[16'h30C7] <= 0;
        weight_mem[16'h30C8] <= 0;
        weight_mem[16'h30C9] <= 0;
        weight_mem[16'h30CA] <= 0;
        weight_mem[16'h30CB] <= 0;
        weight_mem[16'h30CC] <= 0;
        weight_mem[16'h30CD] <= 0;
        weight_mem[16'h30CE] <= 0;
        weight_mem[16'h30CF] <= 0;
        weight_mem[16'h30D0] <= 0;
        weight_mem[16'h30D1] <= 0;
        weight_mem[16'h30D2] <= 0;
        weight_mem[16'h30D3] <= 0;
        weight_mem[16'h30D4] <= 0;
        weight_mem[16'h30D5] <= 0;
        weight_mem[16'h30D6] <= 0;
        weight_mem[16'h30D7] <= 0;
        weight_mem[16'h30D8] <= 0;
        weight_mem[16'h30D9] <= 0;
        weight_mem[16'h30DA] <= 0;
        weight_mem[16'h30DB] <= 0;
        weight_mem[16'h30DC] <= 0;
        weight_mem[16'h30DD] <= 0;
        weight_mem[16'h30DE] <= 0;
        weight_mem[16'h30DF] <= 0;
        weight_mem[16'h30E0] <= 0;
        weight_mem[16'h30E1] <= 0;
        weight_mem[16'h30E2] <= 0;
        weight_mem[16'h30E3] <= 0;
        weight_mem[16'h30E4] <= 0;
        weight_mem[16'h30E5] <= 0;
        weight_mem[16'h30E6] <= 0;
        weight_mem[16'h30E7] <= 0;
        weight_mem[16'h30E8] <= 0;
        weight_mem[16'h30E9] <= 0;
        weight_mem[16'h30EA] <= 0;
        weight_mem[16'h30EB] <= 0;
        weight_mem[16'h30EC] <= 0;
        weight_mem[16'h30ED] <= 0;
        weight_mem[16'h30EE] <= 0;
        weight_mem[16'h30EF] <= 0;
        weight_mem[16'h30F0] <= 0;
        weight_mem[16'h30F1] <= 0;
        weight_mem[16'h30F2] <= 0;
        weight_mem[16'h30F3] <= 0;
        weight_mem[16'h30F4] <= 0;
        weight_mem[16'h30F5] <= 0;
        weight_mem[16'h30F6] <= 0;
        weight_mem[16'h30F7] <= 0;
        weight_mem[16'h30F8] <= 0;
        weight_mem[16'h30F9] <= 0;
        weight_mem[16'h30FA] <= 0;
        weight_mem[16'h30FB] <= 0;
        weight_mem[16'h30FC] <= 0;
        weight_mem[16'h30FD] <= 0;
        weight_mem[16'h30FE] <= 0;
        weight_mem[16'h30FF] <= 0;
        weight_mem[16'h3100] <= 0;
        weight_mem[16'h3101] <= 0;
        weight_mem[16'h3102] <= 0;
        weight_mem[16'h3103] <= 0;
        weight_mem[16'h3104] <= 0;
        weight_mem[16'h3105] <= 0;
        weight_mem[16'h3106] <= 0;
        weight_mem[16'h3107] <= 0;
        weight_mem[16'h3108] <= 0;
        weight_mem[16'h3109] <= 0;
        weight_mem[16'h310A] <= 0;
        weight_mem[16'h310B] <= 0;
        weight_mem[16'h310C] <= 0;
        weight_mem[16'h310D] <= 0;
        weight_mem[16'h310E] <= 0;
        weight_mem[16'h310F] <= 0;
        weight_mem[16'h3110] <= 0;
        weight_mem[16'h3111] <= 0;
        weight_mem[16'h3112] <= 0;
        weight_mem[16'h3113] <= 0;
        weight_mem[16'h3114] <= 0;
        weight_mem[16'h3115] <= 0;
        weight_mem[16'h3116] <= 0;
        weight_mem[16'h3117] <= 0;
        weight_mem[16'h3118] <= 0;
        weight_mem[16'h3119] <= 0;
        weight_mem[16'h311A] <= 0;
        weight_mem[16'h311B] <= 0;
        weight_mem[16'h311C] <= 0;
        weight_mem[16'h311D] <= 0;
        weight_mem[16'h311E] <= 0;
        weight_mem[16'h311F] <= 0;
        weight_mem[16'h3120] <= 0;
        weight_mem[16'h3121] <= 0;
        weight_mem[16'h3122] <= 0;
        weight_mem[16'h3123] <= 0;
        weight_mem[16'h3124] <= 0;
        weight_mem[16'h3125] <= 0;
        weight_mem[16'h3126] <= 0;
        weight_mem[16'h3127] <= 0;
        weight_mem[16'h3128] <= 0;
        weight_mem[16'h3129] <= 0;
        weight_mem[16'h312A] <= 0;
        weight_mem[16'h312B] <= 0;
        weight_mem[16'h312C] <= 0;
        weight_mem[16'h312D] <= 0;
        weight_mem[16'h312E] <= 0;
        weight_mem[16'h312F] <= 0;
        weight_mem[16'h3130] <= 0;
        weight_mem[16'h3131] <= 0;
        weight_mem[16'h3132] <= 0;
        weight_mem[16'h3133] <= 0;
        weight_mem[16'h3134] <= 0;
        weight_mem[16'h3135] <= 0;
        weight_mem[16'h3136] <= 0;
        weight_mem[16'h3137] <= 0;
        weight_mem[16'h3138] <= 0;
        weight_mem[16'h3139] <= 0;
        weight_mem[16'h313A] <= 0;
        weight_mem[16'h313B] <= 0;
        weight_mem[16'h313C] <= 0;
        weight_mem[16'h313D] <= 0;
        weight_mem[16'h313E] <= 0;
        weight_mem[16'h313F] <= 0;
        weight_mem[16'h3140] <= 0;
        weight_mem[16'h3141] <= 0;
        weight_mem[16'h3142] <= 0;
        weight_mem[16'h3143] <= 0;
        weight_mem[16'h3144] <= 0;
        weight_mem[16'h3145] <= 0;
        weight_mem[16'h3146] <= 0;
        weight_mem[16'h3147] <= 0;
        weight_mem[16'h3148] <= 0;
        weight_mem[16'h3149] <= 0;
        weight_mem[16'h314A] <= 0;
        weight_mem[16'h314B] <= 0;
        weight_mem[16'h314C] <= 0;
        weight_mem[16'h314D] <= 0;
        weight_mem[16'h314E] <= 0;
        weight_mem[16'h314F] <= 0;
        weight_mem[16'h3150] <= 0;
        weight_mem[16'h3151] <= 0;
        weight_mem[16'h3152] <= 0;
        weight_mem[16'h3153] <= 0;
        weight_mem[16'h3154] <= 0;
        weight_mem[16'h3155] <= 0;
        weight_mem[16'h3156] <= 0;
        weight_mem[16'h3157] <= 0;
        weight_mem[16'h3158] <= 0;
        weight_mem[16'h3159] <= 0;
        weight_mem[16'h315A] <= 0;
        weight_mem[16'h315B] <= 0;
        weight_mem[16'h315C] <= 0;
        weight_mem[16'h315D] <= 0;
        weight_mem[16'h315E] <= 0;
        weight_mem[16'h315F] <= 0;
        weight_mem[16'h3160] <= 0;
        weight_mem[16'h3161] <= 0;
        weight_mem[16'h3162] <= 0;
        weight_mem[16'h3163] <= 0;
        weight_mem[16'h3164] <= 0;
        weight_mem[16'h3165] <= 0;
        weight_mem[16'h3166] <= 0;
        weight_mem[16'h3167] <= 0;
        weight_mem[16'h3168] <= 0;
        weight_mem[16'h3169] <= 0;
        weight_mem[16'h316A] <= 0;
        weight_mem[16'h316B] <= 0;
        weight_mem[16'h316C] <= 0;
        weight_mem[16'h316D] <= 0;
        weight_mem[16'h316E] <= 0;
        weight_mem[16'h316F] <= 0;
        weight_mem[16'h3170] <= 0;
        weight_mem[16'h3171] <= 0;
        weight_mem[16'h3172] <= 0;
        weight_mem[16'h3173] <= 0;
        weight_mem[16'h3174] <= 0;
        weight_mem[16'h3175] <= 0;
        weight_mem[16'h3176] <= 0;
        weight_mem[16'h3177] <= 0;
        weight_mem[16'h3178] <= 0;
        weight_mem[16'h3179] <= 0;
        weight_mem[16'h317A] <= 0;
        weight_mem[16'h317B] <= 0;
        weight_mem[16'h317C] <= 0;
        weight_mem[16'h317D] <= 0;
        weight_mem[16'h317E] <= 0;
        weight_mem[16'h317F] <= 0;
        weight_mem[16'h3180] <= 0;
        weight_mem[16'h3181] <= 0;
        weight_mem[16'h3182] <= 0;
        weight_mem[16'h3183] <= 0;
        weight_mem[16'h3184] <= 0;
        weight_mem[16'h3185] <= 0;
        weight_mem[16'h3186] <= 0;
        weight_mem[16'h3187] <= 0;
        weight_mem[16'h3188] <= 0;
        weight_mem[16'h3189] <= 0;
        weight_mem[16'h318A] <= 0;
        weight_mem[16'h318B] <= 0;
        weight_mem[16'h318C] <= 0;
        weight_mem[16'h318D] <= 0;
        weight_mem[16'h318E] <= 0;
        weight_mem[16'h318F] <= 0;
        weight_mem[16'h3190] <= 0;
        weight_mem[16'h3191] <= 0;
        weight_mem[16'h3192] <= 0;
        weight_mem[16'h3193] <= 0;
        weight_mem[16'h3194] <= 0;
        weight_mem[16'h3195] <= 0;
        weight_mem[16'h3196] <= 0;
        weight_mem[16'h3197] <= 0;
        weight_mem[16'h3198] <= 0;
        weight_mem[16'h3199] <= 0;
        weight_mem[16'h319A] <= 0;
        weight_mem[16'h319B] <= 0;
        weight_mem[16'h319C] <= 0;
        weight_mem[16'h319D] <= 0;
        weight_mem[16'h319E] <= 0;
        weight_mem[16'h319F] <= 0;
        weight_mem[16'h31A0] <= 0;
        weight_mem[16'h31A1] <= 0;
        weight_mem[16'h31A2] <= 0;
        weight_mem[16'h31A3] <= 0;
        weight_mem[16'h31A4] <= 0;
        weight_mem[16'h31A5] <= 0;
        weight_mem[16'h31A6] <= 0;
        weight_mem[16'h31A7] <= 0;
        weight_mem[16'h31A8] <= 0;
        weight_mem[16'h31A9] <= 0;
        weight_mem[16'h31AA] <= 0;
        weight_mem[16'h31AB] <= 0;
        weight_mem[16'h31AC] <= 0;
        weight_mem[16'h31AD] <= 0;
        weight_mem[16'h31AE] <= 0;
        weight_mem[16'h31AF] <= 0;

        // layer 1 neuron 25
        weight_mem[16'h3200] <= 0;
        weight_mem[16'h3201] <= 0;
        weight_mem[16'h3202] <= 0;
        weight_mem[16'h3203] <= 0;
        weight_mem[16'h3204] <= 0;
        weight_mem[16'h3205] <= 0;
        weight_mem[16'h3206] <= 0;
        weight_mem[16'h3207] <= 0;
        weight_mem[16'h3208] <= 0;
        weight_mem[16'h3209] <= 0;
        weight_mem[16'h320A] <= 0;
        weight_mem[16'h320B] <= 0;
        weight_mem[16'h320C] <= 0;
        weight_mem[16'h320D] <= 0;
        weight_mem[16'h320E] <= 0;
        weight_mem[16'h320F] <= 0;
        weight_mem[16'h3210] <= 0;
        weight_mem[16'h3211] <= 0;
        weight_mem[16'h3212] <= 0;
        weight_mem[16'h3213] <= 0;
        weight_mem[16'h3214] <= 0;
        weight_mem[16'h3215] <= 0;
        weight_mem[16'h3216] <= 0;
        weight_mem[16'h3217] <= 0;
        weight_mem[16'h3218] <= 0;
        weight_mem[16'h3219] <= 0;
        weight_mem[16'h321A] <= 0;
        weight_mem[16'h321B] <= 0;
        weight_mem[16'h321C] <= 0;
        weight_mem[16'h321D] <= 0;
        weight_mem[16'h321E] <= 0;
        weight_mem[16'h321F] <= 0;
        weight_mem[16'h3220] <= 0;
        weight_mem[16'h3221] <= 0;
        weight_mem[16'h3222] <= 0;
        weight_mem[16'h3223] <= 0;
        weight_mem[16'h3224] <= 0;
        weight_mem[16'h3225] <= 0;
        weight_mem[16'h3226] <= 0;
        weight_mem[16'h3227] <= 0;
        weight_mem[16'h3228] <= 0;
        weight_mem[16'h3229] <= 0;
        weight_mem[16'h322A] <= 0;
        weight_mem[16'h322B] <= 0;
        weight_mem[16'h322C] <= 0;
        weight_mem[16'h322D] <= 0;
        weight_mem[16'h322E] <= 0;
        weight_mem[16'h322F] <= 0;
        weight_mem[16'h3230] <= 0;
        weight_mem[16'h3231] <= 0;
        weight_mem[16'h3232] <= 0;
        weight_mem[16'h3233] <= 0;
        weight_mem[16'h3234] <= 0;
        weight_mem[16'h3235] <= 0;
        weight_mem[16'h3236] <= 0;
        weight_mem[16'h3237] <= 0;
        weight_mem[16'h3238] <= 0;
        weight_mem[16'h3239] <= 0;
        weight_mem[16'h323A] <= 0;
        weight_mem[16'h323B] <= 0;
        weight_mem[16'h323C] <= 0;
        weight_mem[16'h323D] <= 0;
        weight_mem[16'h323E] <= 0;
        weight_mem[16'h323F] <= 0;
        weight_mem[16'h3240] <= 0;
        weight_mem[16'h3241] <= 0;
        weight_mem[16'h3242] <= 0;
        weight_mem[16'h3243] <= 0;
        weight_mem[16'h3244] <= 0;
        weight_mem[16'h3245] <= 0;
        weight_mem[16'h3246] <= 0;
        weight_mem[16'h3247] <= 0;
        weight_mem[16'h3248] <= 0;
        weight_mem[16'h3249] <= 0;
        weight_mem[16'h324A] <= 0;
        weight_mem[16'h324B] <= 0;
        weight_mem[16'h324C] <= 0;
        weight_mem[16'h324D] <= 0;
        weight_mem[16'h324E] <= 0;
        weight_mem[16'h324F] <= 0;
        weight_mem[16'h3250] <= 0;
        weight_mem[16'h3251] <= 0;
        weight_mem[16'h3252] <= 0;
        weight_mem[16'h3253] <= 0;
        weight_mem[16'h3254] <= 0;
        weight_mem[16'h3255] <= 0;
        weight_mem[16'h3256] <= 0;
        weight_mem[16'h3257] <= 0;
        weight_mem[16'h3258] <= 0;
        weight_mem[16'h3259] <= 0;
        weight_mem[16'h325A] <= 0;
        weight_mem[16'h325B] <= 0;
        weight_mem[16'h325C] <= 0;
        weight_mem[16'h325D] <= 0;
        weight_mem[16'h325E] <= 0;
        weight_mem[16'h325F] <= 0;
        weight_mem[16'h3260] <= 0;
        weight_mem[16'h3261] <= 0;
        weight_mem[16'h3262] <= 0;
        weight_mem[16'h3263] <= 0;
        weight_mem[16'h3264] <= 0;
        weight_mem[16'h3265] <= 0;
        weight_mem[16'h3266] <= 0;
        weight_mem[16'h3267] <= 0;
        weight_mem[16'h3268] <= 0;
        weight_mem[16'h3269] <= 0;
        weight_mem[16'h326A] <= 0;
        weight_mem[16'h326B] <= 0;
        weight_mem[16'h326C] <= 0;
        weight_mem[16'h326D] <= 0;
        weight_mem[16'h326E] <= 0;
        weight_mem[16'h326F] <= 0;
        weight_mem[16'h3270] <= 0;
        weight_mem[16'h3271] <= 0;
        weight_mem[16'h3272] <= 0;
        weight_mem[16'h3273] <= 0;
        weight_mem[16'h3274] <= 0;
        weight_mem[16'h3275] <= 0;
        weight_mem[16'h3276] <= 0;
        weight_mem[16'h3277] <= 0;
        weight_mem[16'h3278] <= 0;
        weight_mem[16'h3279] <= 0;
        weight_mem[16'h327A] <= 0;
        weight_mem[16'h327B] <= 0;
        weight_mem[16'h327C] <= 0;
        weight_mem[16'h327D] <= 0;
        weight_mem[16'h327E] <= 0;
        weight_mem[16'h327F] <= 0;
        weight_mem[16'h3280] <= 0;
        weight_mem[16'h3281] <= 0;
        weight_mem[16'h3282] <= 0;
        weight_mem[16'h3283] <= 0;
        weight_mem[16'h3284] <= 0;
        weight_mem[16'h3285] <= 0;
        weight_mem[16'h3286] <= 0;
        weight_mem[16'h3287] <= 0;
        weight_mem[16'h3288] <= 0;
        weight_mem[16'h3289] <= 0;
        weight_mem[16'h328A] <= 0;
        weight_mem[16'h328B] <= 0;
        weight_mem[16'h328C] <= 0;
        weight_mem[16'h328D] <= 0;
        weight_mem[16'h328E] <= 0;
        weight_mem[16'h328F] <= 0;
        weight_mem[16'h3290] <= 0;
        weight_mem[16'h3291] <= 0;
        weight_mem[16'h3292] <= 0;
        weight_mem[16'h3293] <= 0;
        weight_mem[16'h3294] <= 0;
        weight_mem[16'h3295] <= 0;
        weight_mem[16'h3296] <= 0;
        weight_mem[16'h3297] <= 0;
        weight_mem[16'h3298] <= 0;
        weight_mem[16'h3299] <= 0;
        weight_mem[16'h329A] <= 0;
        weight_mem[16'h329B] <= 0;
        weight_mem[16'h329C] <= 0;
        weight_mem[16'h329D] <= 0;
        weight_mem[16'h329E] <= 0;
        weight_mem[16'h329F] <= 0;
        weight_mem[16'h32A0] <= 0;
        weight_mem[16'h32A1] <= 0;
        weight_mem[16'h32A2] <= 0;
        weight_mem[16'h32A3] <= 0;
        weight_mem[16'h32A4] <= 0;
        weight_mem[16'h32A5] <= 0;
        weight_mem[16'h32A6] <= 0;
        weight_mem[16'h32A7] <= 0;
        weight_mem[16'h32A8] <= 0;
        weight_mem[16'h32A9] <= 0;
        weight_mem[16'h32AA] <= 0;
        weight_mem[16'h32AB] <= 0;
        weight_mem[16'h32AC] <= 0;
        weight_mem[16'h32AD] <= 0;
        weight_mem[16'h32AE] <= 0;
        weight_mem[16'h32AF] <= 0;
        weight_mem[16'h32B0] <= 0;
        weight_mem[16'h32B1] <= 0;
        weight_mem[16'h32B2] <= 0;
        weight_mem[16'h32B3] <= 0;
        weight_mem[16'h32B4] <= 0;
        weight_mem[16'h32B5] <= 0;
        weight_mem[16'h32B6] <= 0;
        weight_mem[16'h32B7] <= 0;
        weight_mem[16'h32B8] <= 0;
        weight_mem[16'h32B9] <= 0;
        weight_mem[16'h32BA] <= 0;
        weight_mem[16'h32BB] <= 0;
        weight_mem[16'h32BC] <= 0;
        weight_mem[16'h32BD] <= 0;
        weight_mem[16'h32BE] <= 0;
        weight_mem[16'h32BF] <= 0;
        weight_mem[16'h32C0] <= 0;
        weight_mem[16'h32C1] <= 0;
        weight_mem[16'h32C2] <= 0;
        weight_mem[16'h32C3] <= 0;
        weight_mem[16'h32C4] <= 0;
        weight_mem[16'h32C5] <= 0;
        weight_mem[16'h32C6] <= 0;
        weight_mem[16'h32C7] <= 0;
        weight_mem[16'h32C8] <= 0;
        weight_mem[16'h32C9] <= 0;
        weight_mem[16'h32CA] <= 0;
        weight_mem[16'h32CB] <= 0;
        weight_mem[16'h32CC] <= 0;
        weight_mem[16'h32CD] <= 0;
        weight_mem[16'h32CE] <= 0;
        weight_mem[16'h32CF] <= 0;
        weight_mem[16'h32D0] <= 0;
        weight_mem[16'h32D1] <= 0;
        weight_mem[16'h32D2] <= 0;
        weight_mem[16'h32D3] <= 0;
        weight_mem[16'h32D4] <= 0;
        weight_mem[16'h32D5] <= 0;
        weight_mem[16'h32D6] <= 0;
        weight_mem[16'h32D7] <= 0;
        weight_mem[16'h32D8] <= 0;
        weight_mem[16'h32D9] <= 0;
        weight_mem[16'h32DA] <= 0;
        weight_mem[16'h32DB] <= 0;
        weight_mem[16'h32DC] <= 0;
        weight_mem[16'h32DD] <= 0;
        weight_mem[16'h32DE] <= 0;
        weight_mem[16'h32DF] <= 0;
        weight_mem[16'h32E0] <= 0;
        weight_mem[16'h32E1] <= 0;
        weight_mem[16'h32E2] <= 0;
        weight_mem[16'h32E3] <= 0;
        weight_mem[16'h32E4] <= 0;
        weight_mem[16'h32E5] <= 0;
        weight_mem[16'h32E6] <= 0;
        weight_mem[16'h32E7] <= 0;
        weight_mem[16'h32E8] <= 0;
        weight_mem[16'h32E9] <= 0;
        weight_mem[16'h32EA] <= 0;
        weight_mem[16'h32EB] <= 0;
        weight_mem[16'h32EC] <= 0;
        weight_mem[16'h32ED] <= 0;
        weight_mem[16'h32EE] <= 0;
        weight_mem[16'h32EF] <= 0;
        weight_mem[16'h32F0] <= 0;
        weight_mem[16'h32F1] <= 0;
        weight_mem[16'h32F2] <= 0;
        weight_mem[16'h32F3] <= 0;
        weight_mem[16'h32F4] <= 0;
        weight_mem[16'h32F5] <= 0;
        weight_mem[16'h32F6] <= 0;
        weight_mem[16'h32F7] <= 0;
        weight_mem[16'h32F8] <= 0;
        weight_mem[16'h32F9] <= 0;
        weight_mem[16'h32FA] <= 0;
        weight_mem[16'h32FB] <= 0;
        weight_mem[16'h32FC] <= 0;
        weight_mem[16'h32FD] <= 0;
        weight_mem[16'h32FE] <= 0;
        weight_mem[16'h32FF] <= 0;
        weight_mem[16'h3300] <= 0;
        weight_mem[16'h3301] <= 0;
        weight_mem[16'h3302] <= 0;
        weight_mem[16'h3303] <= 0;
        weight_mem[16'h3304] <= 0;
        weight_mem[16'h3305] <= 0;
        weight_mem[16'h3306] <= 0;
        weight_mem[16'h3307] <= 0;
        weight_mem[16'h3308] <= 0;
        weight_mem[16'h3309] <= 0;
        weight_mem[16'h330A] <= 0;
        weight_mem[16'h330B] <= 0;
        weight_mem[16'h330C] <= 0;
        weight_mem[16'h330D] <= 0;
        weight_mem[16'h330E] <= 0;
        weight_mem[16'h330F] <= 0;
        weight_mem[16'h3310] <= 0;
        weight_mem[16'h3311] <= 0;
        weight_mem[16'h3312] <= 0;
        weight_mem[16'h3313] <= 0;
        weight_mem[16'h3314] <= 0;
        weight_mem[16'h3315] <= 0;
        weight_mem[16'h3316] <= 0;
        weight_mem[16'h3317] <= 0;
        weight_mem[16'h3318] <= 0;
        weight_mem[16'h3319] <= 0;
        weight_mem[16'h331A] <= 0;
        weight_mem[16'h331B] <= 0;
        weight_mem[16'h331C] <= 0;
        weight_mem[16'h331D] <= 0;
        weight_mem[16'h331E] <= 0;
        weight_mem[16'h331F] <= 0;
        weight_mem[16'h3320] <= 0;
        weight_mem[16'h3321] <= 0;
        weight_mem[16'h3322] <= 0;
        weight_mem[16'h3323] <= 0;
        weight_mem[16'h3324] <= 0;
        weight_mem[16'h3325] <= 0;
        weight_mem[16'h3326] <= 0;
        weight_mem[16'h3327] <= 0;
        weight_mem[16'h3328] <= 0;
        weight_mem[16'h3329] <= 0;
        weight_mem[16'h332A] <= 0;
        weight_mem[16'h332B] <= 0;
        weight_mem[16'h332C] <= 0;
        weight_mem[16'h332D] <= 0;
        weight_mem[16'h332E] <= 0;
        weight_mem[16'h332F] <= 0;
        weight_mem[16'h3330] <= 0;
        weight_mem[16'h3331] <= 0;
        weight_mem[16'h3332] <= 0;
        weight_mem[16'h3333] <= 0;
        weight_mem[16'h3334] <= 0;
        weight_mem[16'h3335] <= 0;
        weight_mem[16'h3336] <= 0;
        weight_mem[16'h3337] <= 0;
        weight_mem[16'h3338] <= 0;
        weight_mem[16'h3339] <= 0;
        weight_mem[16'h333A] <= 0;
        weight_mem[16'h333B] <= 0;
        weight_mem[16'h333C] <= 0;
        weight_mem[16'h333D] <= 0;
        weight_mem[16'h333E] <= 0;
        weight_mem[16'h333F] <= 0;
        weight_mem[16'h3340] <= 0;
        weight_mem[16'h3341] <= 0;
        weight_mem[16'h3342] <= 0;
        weight_mem[16'h3343] <= 0;
        weight_mem[16'h3344] <= 0;
        weight_mem[16'h3345] <= 0;
        weight_mem[16'h3346] <= 0;
        weight_mem[16'h3347] <= 0;
        weight_mem[16'h3348] <= 0;
        weight_mem[16'h3349] <= 0;
        weight_mem[16'h334A] <= 0;
        weight_mem[16'h334B] <= 0;
        weight_mem[16'h334C] <= 0;
        weight_mem[16'h334D] <= 0;
        weight_mem[16'h334E] <= 0;
        weight_mem[16'h334F] <= 0;
        weight_mem[16'h3350] <= 0;
        weight_mem[16'h3351] <= 0;
        weight_mem[16'h3352] <= 0;
        weight_mem[16'h3353] <= 0;
        weight_mem[16'h3354] <= 0;
        weight_mem[16'h3355] <= 0;
        weight_mem[16'h3356] <= 0;
        weight_mem[16'h3357] <= 0;
        weight_mem[16'h3358] <= 0;
        weight_mem[16'h3359] <= 0;
        weight_mem[16'h335A] <= 0;
        weight_mem[16'h335B] <= 0;
        weight_mem[16'h335C] <= 0;
        weight_mem[16'h335D] <= 0;
        weight_mem[16'h335E] <= 0;
        weight_mem[16'h335F] <= 0;
        weight_mem[16'h3360] <= 0;
        weight_mem[16'h3361] <= 0;
        weight_mem[16'h3362] <= 0;
        weight_mem[16'h3363] <= 0;
        weight_mem[16'h3364] <= 0;
        weight_mem[16'h3365] <= 0;
        weight_mem[16'h3366] <= 0;
        weight_mem[16'h3367] <= 0;
        weight_mem[16'h3368] <= 0;
        weight_mem[16'h3369] <= 0;
        weight_mem[16'h336A] <= 0;
        weight_mem[16'h336B] <= 0;
        weight_mem[16'h336C] <= 0;
        weight_mem[16'h336D] <= 0;
        weight_mem[16'h336E] <= 0;
        weight_mem[16'h336F] <= 0;
        weight_mem[16'h3370] <= 0;
        weight_mem[16'h3371] <= 0;
        weight_mem[16'h3372] <= 0;
        weight_mem[16'h3373] <= 0;
        weight_mem[16'h3374] <= 0;
        weight_mem[16'h3375] <= 0;
        weight_mem[16'h3376] <= 0;
        weight_mem[16'h3377] <= 0;
        weight_mem[16'h3378] <= 0;
        weight_mem[16'h3379] <= 0;
        weight_mem[16'h337A] <= 0;
        weight_mem[16'h337B] <= 0;
        weight_mem[16'h337C] <= 0;
        weight_mem[16'h337D] <= 0;
        weight_mem[16'h337E] <= 0;
        weight_mem[16'h337F] <= 0;
        weight_mem[16'h3380] <= 0;
        weight_mem[16'h3381] <= 0;
        weight_mem[16'h3382] <= 0;
        weight_mem[16'h3383] <= 0;
        weight_mem[16'h3384] <= 0;
        weight_mem[16'h3385] <= 0;
        weight_mem[16'h3386] <= 0;
        weight_mem[16'h3387] <= 0;
        weight_mem[16'h3388] <= 0;
        weight_mem[16'h3389] <= 0;
        weight_mem[16'h338A] <= 0;
        weight_mem[16'h338B] <= 0;
        weight_mem[16'h338C] <= 0;
        weight_mem[16'h338D] <= 0;
        weight_mem[16'h338E] <= 0;
        weight_mem[16'h338F] <= 0;
        weight_mem[16'h3390] <= 0;
        weight_mem[16'h3391] <= 0;
        weight_mem[16'h3392] <= 0;
        weight_mem[16'h3393] <= 0;
        weight_mem[16'h3394] <= 0;
        weight_mem[16'h3395] <= 0;
        weight_mem[16'h3396] <= 0;
        weight_mem[16'h3397] <= 0;
        weight_mem[16'h3398] <= 0;
        weight_mem[16'h3399] <= 0;
        weight_mem[16'h339A] <= 0;
        weight_mem[16'h339B] <= 0;
        weight_mem[16'h339C] <= 0;
        weight_mem[16'h339D] <= 0;
        weight_mem[16'h339E] <= 0;
        weight_mem[16'h339F] <= 0;
        weight_mem[16'h33A0] <= 0;
        weight_mem[16'h33A1] <= 0;
        weight_mem[16'h33A2] <= 0;
        weight_mem[16'h33A3] <= 0;
        weight_mem[16'h33A4] <= 0;
        weight_mem[16'h33A5] <= 0;
        weight_mem[16'h33A6] <= 0;
        weight_mem[16'h33A7] <= 0;
        weight_mem[16'h33A8] <= 0;
        weight_mem[16'h33A9] <= 0;
        weight_mem[16'h33AA] <= 0;
        weight_mem[16'h33AB] <= 0;
        weight_mem[16'h33AC] <= 0;
        weight_mem[16'h33AD] <= 0;
        weight_mem[16'h33AE] <= 0;
        weight_mem[16'h33AF] <= 0;

        // layer 1 neuron 26
        weight_mem[16'h3400] <= 0;
        weight_mem[16'h3401] <= 0;
        weight_mem[16'h3402] <= 0;
        weight_mem[16'h3403] <= 0;
        weight_mem[16'h3404] <= 0;
        weight_mem[16'h3405] <= 0;
        weight_mem[16'h3406] <= 0;
        weight_mem[16'h3407] <= 0;
        weight_mem[16'h3408] <= 0;
        weight_mem[16'h3409] <= 0;
        weight_mem[16'h340A] <= 0;
        weight_mem[16'h340B] <= 0;
        weight_mem[16'h340C] <= 0;
        weight_mem[16'h340D] <= 0;
        weight_mem[16'h340E] <= 0;
        weight_mem[16'h340F] <= 0;
        weight_mem[16'h3410] <= 0;
        weight_mem[16'h3411] <= 0;
        weight_mem[16'h3412] <= 0;
        weight_mem[16'h3413] <= 0;
        weight_mem[16'h3414] <= 0;
        weight_mem[16'h3415] <= 0;
        weight_mem[16'h3416] <= 0;
        weight_mem[16'h3417] <= 0;
        weight_mem[16'h3418] <= 0;
        weight_mem[16'h3419] <= 0;
        weight_mem[16'h341A] <= 0;
        weight_mem[16'h341B] <= 0;
        weight_mem[16'h341C] <= 0;
        weight_mem[16'h341D] <= 0;
        weight_mem[16'h341E] <= 0;
        weight_mem[16'h341F] <= 0;
        weight_mem[16'h3420] <= 0;
        weight_mem[16'h3421] <= 0;
        weight_mem[16'h3422] <= 0;
        weight_mem[16'h3423] <= 0;
        weight_mem[16'h3424] <= 0;
        weight_mem[16'h3425] <= 0;
        weight_mem[16'h3426] <= 0;
        weight_mem[16'h3427] <= 0;
        weight_mem[16'h3428] <= 0;
        weight_mem[16'h3429] <= 0;
        weight_mem[16'h342A] <= 0;
        weight_mem[16'h342B] <= 0;
        weight_mem[16'h342C] <= 0;
        weight_mem[16'h342D] <= 0;
        weight_mem[16'h342E] <= 0;
        weight_mem[16'h342F] <= 0;
        weight_mem[16'h3430] <= 0;
        weight_mem[16'h3431] <= 0;
        weight_mem[16'h3432] <= 0;
        weight_mem[16'h3433] <= 0;
        weight_mem[16'h3434] <= 0;
        weight_mem[16'h3435] <= 0;
        weight_mem[16'h3436] <= 0;
        weight_mem[16'h3437] <= 0;
        weight_mem[16'h3438] <= 0;
        weight_mem[16'h3439] <= 0;
        weight_mem[16'h343A] <= 0;
        weight_mem[16'h343B] <= 0;
        weight_mem[16'h343C] <= 0;
        weight_mem[16'h343D] <= 0;
        weight_mem[16'h343E] <= 0;
        weight_mem[16'h343F] <= 0;
        weight_mem[16'h3440] <= 0;
        weight_mem[16'h3441] <= 0;
        weight_mem[16'h3442] <= 0;
        weight_mem[16'h3443] <= 0;
        weight_mem[16'h3444] <= 0;
        weight_mem[16'h3445] <= 0;
        weight_mem[16'h3446] <= 0;
        weight_mem[16'h3447] <= 0;
        weight_mem[16'h3448] <= 0;
        weight_mem[16'h3449] <= 0;
        weight_mem[16'h344A] <= 0;
        weight_mem[16'h344B] <= 0;
        weight_mem[16'h344C] <= 0;
        weight_mem[16'h344D] <= 0;
        weight_mem[16'h344E] <= 0;
        weight_mem[16'h344F] <= 0;
        weight_mem[16'h3450] <= 0;
        weight_mem[16'h3451] <= 0;
        weight_mem[16'h3452] <= 0;
        weight_mem[16'h3453] <= 0;
        weight_mem[16'h3454] <= 0;
        weight_mem[16'h3455] <= 0;
        weight_mem[16'h3456] <= 0;
        weight_mem[16'h3457] <= 0;
        weight_mem[16'h3458] <= 0;
        weight_mem[16'h3459] <= 0;
        weight_mem[16'h345A] <= 0;
        weight_mem[16'h345B] <= 0;
        weight_mem[16'h345C] <= 0;
        weight_mem[16'h345D] <= 0;
        weight_mem[16'h345E] <= 0;
        weight_mem[16'h345F] <= 0;
        weight_mem[16'h3460] <= 0;
        weight_mem[16'h3461] <= 0;
        weight_mem[16'h3462] <= 0;
        weight_mem[16'h3463] <= 0;
        weight_mem[16'h3464] <= 0;
        weight_mem[16'h3465] <= 0;
        weight_mem[16'h3466] <= 0;
        weight_mem[16'h3467] <= 0;
        weight_mem[16'h3468] <= 0;
        weight_mem[16'h3469] <= 0;
        weight_mem[16'h346A] <= 0;
        weight_mem[16'h346B] <= 0;
        weight_mem[16'h346C] <= 0;
        weight_mem[16'h346D] <= 0;
        weight_mem[16'h346E] <= 0;
        weight_mem[16'h346F] <= 0;
        weight_mem[16'h3470] <= 0;
        weight_mem[16'h3471] <= 0;
        weight_mem[16'h3472] <= 0;
        weight_mem[16'h3473] <= 0;
        weight_mem[16'h3474] <= 0;
        weight_mem[16'h3475] <= 0;
        weight_mem[16'h3476] <= 0;
        weight_mem[16'h3477] <= 0;
        weight_mem[16'h3478] <= 0;
        weight_mem[16'h3479] <= 0;
        weight_mem[16'h347A] <= 0;
        weight_mem[16'h347B] <= 0;
        weight_mem[16'h347C] <= 0;
        weight_mem[16'h347D] <= 0;
        weight_mem[16'h347E] <= 0;
        weight_mem[16'h347F] <= 0;
        weight_mem[16'h3480] <= 0;
        weight_mem[16'h3481] <= 0;
        weight_mem[16'h3482] <= 0;
        weight_mem[16'h3483] <= 0;
        weight_mem[16'h3484] <= 0;
        weight_mem[16'h3485] <= 0;
        weight_mem[16'h3486] <= 0;
        weight_mem[16'h3487] <= 0;
        weight_mem[16'h3488] <= 0;
        weight_mem[16'h3489] <= 0;
        weight_mem[16'h348A] <= 0;
        weight_mem[16'h348B] <= 0;
        weight_mem[16'h348C] <= 0;
        weight_mem[16'h348D] <= 0;
        weight_mem[16'h348E] <= 0;
        weight_mem[16'h348F] <= 0;
        weight_mem[16'h3490] <= 0;
        weight_mem[16'h3491] <= 0;
        weight_mem[16'h3492] <= 0;
        weight_mem[16'h3493] <= 0;
        weight_mem[16'h3494] <= 0;
        weight_mem[16'h3495] <= 0;
        weight_mem[16'h3496] <= 0;
        weight_mem[16'h3497] <= 0;
        weight_mem[16'h3498] <= 0;
        weight_mem[16'h3499] <= 0;
        weight_mem[16'h349A] <= 0;
        weight_mem[16'h349B] <= 0;
        weight_mem[16'h349C] <= 0;
        weight_mem[16'h349D] <= 0;
        weight_mem[16'h349E] <= 0;
        weight_mem[16'h349F] <= 0;
        weight_mem[16'h34A0] <= 0;
        weight_mem[16'h34A1] <= 0;
        weight_mem[16'h34A2] <= 0;
        weight_mem[16'h34A3] <= 0;
        weight_mem[16'h34A4] <= 0;
        weight_mem[16'h34A5] <= 0;
        weight_mem[16'h34A6] <= 0;
        weight_mem[16'h34A7] <= 0;
        weight_mem[16'h34A8] <= 0;
        weight_mem[16'h34A9] <= 0;
        weight_mem[16'h34AA] <= 0;
        weight_mem[16'h34AB] <= 0;
        weight_mem[16'h34AC] <= 0;
        weight_mem[16'h34AD] <= 0;
        weight_mem[16'h34AE] <= 0;
        weight_mem[16'h34AF] <= 0;
        weight_mem[16'h34B0] <= 0;
        weight_mem[16'h34B1] <= 0;
        weight_mem[16'h34B2] <= 0;
        weight_mem[16'h34B3] <= 0;
        weight_mem[16'h34B4] <= 0;
        weight_mem[16'h34B5] <= 0;
        weight_mem[16'h34B6] <= 0;
        weight_mem[16'h34B7] <= 0;
        weight_mem[16'h34B8] <= 0;
        weight_mem[16'h34B9] <= 0;
        weight_mem[16'h34BA] <= 0;
        weight_mem[16'h34BB] <= 0;
        weight_mem[16'h34BC] <= 0;
        weight_mem[16'h34BD] <= 0;
        weight_mem[16'h34BE] <= 0;
        weight_mem[16'h34BF] <= 0;
        weight_mem[16'h34C0] <= 0;
        weight_mem[16'h34C1] <= 0;
        weight_mem[16'h34C2] <= 0;
        weight_mem[16'h34C3] <= 0;
        weight_mem[16'h34C4] <= 0;
        weight_mem[16'h34C5] <= 0;
        weight_mem[16'h34C6] <= 0;
        weight_mem[16'h34C7] <= 0;
        weight_mem[16'h34C8] <= 0;
        weight_mem[16'h34C9] <= 0;
        weight_mem[16'h34CA] <= 0;
        weight_mem[16'h34CB] <= 0;
        weight_mem[16'h34CC] <= 0;
        weight_mem[16'h34CD] <= 0;
        weight_mem[16'h34CE] <= 0;
        weight_mem[16'h34CF] <= 0;
        weight_mem[16'h34D0] <= 0;
        weight_mem[16'h34D1] <= 0;
        weight_mem[16'h34D2] <= 0;
        weight_mem[16'h34D3] <= 0;
        weight_mem[16'h34D4] <= 0;
        weight_mem[16'h34D5] <= 0;
        weight_mem[16'h34D6] <= 0;
        weight_mem[16'h34D7] <= 0;
        weight_mem[16'h34D8] <= 0;
        weight_mem[16'h34D9] <= 0;
        weight_mem[16'h34DA] <= 0;
        weight_mem[16'h34DB] <= 0;
        weight_mem[16'h34DC] <= 0;
        weight_mem[16'h34DD] <= 0;
        weight_mem[16'h34DE] <= 0;
        weight_mem[16'h34DF] <= 0;
        weight_mem[16'h34E0] <= 0;
        weight_mem[16'h34E1] <= 0;
        weight_mem[16'h34E2] <= 0;
        weight_mem[16'h34E3] <= 0;
        weight_mem[16'h34E4] <= 0;
        weight_mem[16'h34E5] <= 0;
        weight_mem[16'h34E6] <= 0;
        weight_mem[16'h34E7] <= 0;
        weight_mem[16'h34E8] <= 0;
        weight_mem[16'h34E9] <= 0;
        weight_mem[16'h34EA] <= 0;
        weight_mem[16'h34EB] <= 0;
        weight_mem[16'h34EC] <= 0;
        weight_mem[16'h34ED] <= 0;
        weight_mem[16'h34EE] <= 0;
        weight_mem[16'h34EF] <= 0;
        weight_mem[16'h34F0] <= 0;
        weight_mem[16'h34F1] <= 0;
        weight_mem[16'h34F2] <= 0;
        weight_mem[16'h34F3] <= 0;
        weight_mem[16'h34F4] <= 0;
        weight_mem[16'h34F5] <= 0;
        weight_mem[16'h34F6] <= 0;
        weight_mem[16'h34F7] <= 0;
        weight_mem[16'h34F8] <= 0;
        weight_mem[16'h34F9] <= 0;
        weight_mem[16'h34FA] <= 0;
        weight_mem[16'h34FB] <= 0;
        weight_mem[16'h34FC] <= 0;
        weight_mem[16'h34FD] <= 0;
        weight_mem[16'h34FE] <= 0;
        weight_mem[16'h34FF] <= 0;
        weight_mem[16'h3500] <= 0;
        weight_mem[16'h3501] <= 0;
        weight_mem[16'h3502] <= 0;
        weight_mem[16'h3503] <= 0;
        weight_mem[16'h3504] <= 0;
        weight_mem[16'h3505] <= 0;
        weight_mem[16'h3506] <= 0;
        weight_mem[16'h3507] <= 0;
        weight_mem[16'h3508] <= 0;
        weight_mem[16'h3509] <= 0;
        weight_mem[16'h350A] <= 0;
        weight_mem[16'h350B] <= 0;
        weight_mem[16'h350C] <= 0;
        weight_mem[16'h350D] <= 0;
        weight_mem[16'h350E] <= 0;
        weight_mem[16'h350F] <= 0;
        weight_mem[16'h3510] <= 0;
        weight_mem[16'h3511] <= 0;
        weight_mem[16'h3512] <= 0;
        weight_mem[16'h3513] <= 0;
        weight_mem[16'h3514] <= 0;
        weight_mem[16'h3515] <= 0;
        weight_mem[16'h3516] <= 0;
        weight_mem[16'h3517] <= 0;
        weight_mem[16'h3518] <= 0;
        weight_mem[16'h3519] <= 0;
        weight_mem[16'h351A] <= 0;
        weight_mem[16'h351B] <= 0;
        weight_mem[16'h351C] <= 0;
        weight_mem[16'h351D] <= 0;
        weight_mem[16'h351E] <= 0;
        weight_mem[16'h351F] <= 0;
        weight_mem[16'h3520] <= 0;
        weight_mem[16'h3521] <= 0;
        weight_mem[16'h3522] <= 0;
        weight_mem[16'h3523] <= 0;
        weight_mem[16'h3524] <= 0;
        weight_mem[16'h3525] <= 0;
        weight_mem[16'h3526] <= 0;
        weight_mem[16'h3527] <= 0;
        weight_mem[16'h3528] <= 0;
        weight_mem[16'h3529] <= 0;
        weight_mem[16'h352A] <= 0;
        weight_mem[16'h352B] <= 0;
        weight_mem[16'h352C] <= 0;
        weight_mem[16'h352D] <= 0;
        weight_mem[16'h352E] <= 0;
        weight_mem[16'h352F] <= 0;
        weight_mem[16'h3530] <= 0;
        weight_mem[16'h3531] <= 0;
        weight_mem[16'h3532] <= 0;
        weight_mem[16'h3533] <= 0;
        weight_mem[16'h3534] <= 0;
        weight_mem[16'h3535] <= 0;
        weight_mem[16'h3536] <= 0;
        weight_mem[16'h3537] <= 0;
        weight_mem[16'h3538] <= 0;
        weight_mem[16'h3539] <= 0;
        weight_mem[16'h353A] <= 0;
        weight_mem[16'h353B] <= 0;
        weight_mem[16'h353C] <= 0;
        weight_mem[16'h353D] <= 0;
        weight_mem[16'h353E] <= 0;
        weight_mem[16'h353F] <= 0;
        weight_mem[16'h3540] <= 0;
        weight_mem[16'h3541] <= 0;
        weight_mem[16'h3542] <= 0;
        weight_mem[16'h3543] <= 0;
        weight_mem[16'h3544] <= 0;
        weight_mem[16'h3545] <= 0;
        weight_mem[16'h3546] <= 0;
        weight_mem[16'h3547] <= 0;
        weight_mem[16'h3548] <= 0;
        weight_mem[16'h3549] <= 0;
        weight_mem[16'h354A] <= 0;
        weight_mem[16'h354B] <= 0;
        weight_mem[16'h354C] <= 0;
        weight_mem[16'h354D] <= 0;
        weight_mem[16'h354E] <= 0;
        weight_mem[16'h354F] <= 0;
        weight_mem[16'h3550] <= 0;
        weight_mem[16'h3551] <= 0;
        weight_mem[16'h3552] <= 0;
        weight_mem[16'h3553] <= 0;
        weight_mem[16'h3554] <= 0;
        weight_mem[16'h3555] <= 0;
        weight_mem[16'h3556] <= 0;
        weight_mem[16'h3557] <= 0;
        weight_mem[16'h3558] <= 0;
        weight_mem[16'h3559] <= 0;
        weight_mem[16'h355A] <= 0;
        weight_mem[16'h355B] <= 0;
        weight_mem[16'h355C] <= 0;
        weight_mem[16'h355D] <= 0;
        weight_mem[16'h355E] <= 0;
        weight_mem[16'h355F] <= 0;
        weight_mem[16'h3560] <= 0;
        weight_mem[16'h3561] <= 0;
        weight_mem[16'h3562] <= 0;
        weight_mem[16'h3563] <= 0;
        weight_mem[16'h3564] <= 0;
        weight_mem[16'h3565] <= 0;
        weight_mem[16'h3566] <= 0;
        weight_mem[16'h3567] <= 0;
        weight_mem[16'h3568] <= 0;
        weight_mem[16'h3569] <= 0;
        weight_mem[16'h356A] <= 0;
        weight_mem[16'h356B] <= 0;
        weight_mem[16'h356C] <= 0;
        weight_mem[16'h356D] <= 0;
        weight_mem[16'h356E] <= 0;
        weight_mem[16'h356F] <= 0;
        weight_mem[16'h3570] <= 0;
        weight_mem[16'h3571] <= 0;
        weight_mem[16'h3572] <= 0;
        weight_mem[16'h3573] <= 0;
        weight_mem[16'h3574] <= 0;
        weight_mem[16'h3575] <= 0;
        weight_mem[16'h3576] <= 0;
        weight_mem[16'h3577] <= 0;
        weight_mem[16'h3578] <= 0;
        weight_mem[16'h3579] <= 0;
        weight_mem[16'h357A] <= 0;
        weight_mem[16'h357B] <= 0;
        weight_mem[16'h357C] <= 0;
        weight_mem[16'h357D] <= 0;
        weight_mem[16'h357E] <= 0;
        weight_mem[16'h357F] <= 0;
        weight_mem[16'h3580] <= 0;
        weight_mem[16'h3581] <= 0;
        weight_mem[16'h3582] <= 0;
        weight_mem[16'h3583] <= 0;
        weight_mem[16'h3584] <= 0;
        weight_mem[16'h3585] <= 0;
        weight_mem[16'h3586] <= 0;
        weight_mem[16'h3587] <= 0;
        weight_mem[16'h3588] <= 0;
        weight_mem[16'h3589] <= 0;
        weight_mem[16'h358A] <= 0;
        weight_mem[16'h358B] <= 0;
        weight_mem[16'h358C] <= 0;
        weight_mem[16'h358D] <= 0;
        weight_mem[16'h358E] <= 0;
        weight_mem[16'h358F] <= 0;
        weight_mem[16'h3590] <= 0;
        weight_mem[16'h3591] <= 0;
        weight_mem[16'h3592] <= 0;
        weight_mem[16'h3593] <= 0;
        weight_mem[16'h3594] <= 0;
        weight_mem[16'h3595] <= 0;
        weight_mem[16'h3596] <= 0;
        weight_mem[16'h3597] <= 0;
        weight_mem[16'h3598] <= 0;
        weight_mem[16'h3599] <= 0;
        weight_mem[16'h359A] <= 0;
        weight_mem[16'h359B] <= 0;
        weight_mem[16'h359C] <= 0;
        weight_mem[16'h359D] <= 0;
        weight_mem[16'h359E] <= 0;
        weight_mem[16'h359F] <= 0;
        weight_mem[16'h35A0] <= 0;
        weight_mem[16'h35A1] <= 0;
        weight_mem[16'h35A2] <= 0;
        weight_mem[16'h35A3] <= 0;
        weight_mem[16'h35A4] <= 0;
        weight_mem[16'h35A5] <= 0;
        weight_mem[16'h35A6] <= 0;
        weight_mem[16'h35A7] <= 0;
        weight_mem[16'h35A8] <= 0;
        weight_mem[16'h35A9] <= 0;
        weight_mem[16'h35AA] <= 0;
        weight_mem[16'h35AB] <= 0;
        weight_mem[16'h35AC] <= 0;
        weight_mem[16'h35AD] <= 0;
        weight_mem[16'h35AE] <= 0;
        weight_mem[16'h35AF] <= 0;

        // layer 1 neuron 27
        weight_mem[16'h3600] <= 0;
        weight_mem[16'h3601] <= 0;
        weight_mem[16'h3602] <= 0;
        weight_mem[16'h3603] <= 0;
        weight_mem[16'h3604] <= 0;
        weight_mem[16'h3605] <= 0;
        weight_mem[16'h3606] <= 0;
        weight_mem[16'h3607] <= 0;
        weight_mem[16'h3608] <= 0;
        weight_mem[16'h3609] <= 0;
        weight_mem[16'h360A] <= 0;
        weight_mem[16'h360B] <= 0;
        weight_mem[16'h360C] <= 0;
        weight_mem[16'h360D] <= 0;
        weight_mem[16'h360E] <= 0;
        weight_mem[16'h360F] <= 0;
        weight_mem[16'h3610] <= 0;
        weight_mem[16'h3611] <= 0;
        weight_mem[16'h3612] <= 0;
        weight_mem[16'h3613] <= 0;
        weight_mem[16'h3614] <= 0;
        weight_mem[16'h3615] <= 0;
        weight_mem[16'h3616] <= 0;
        weight_mem[16'h3617] <= 0;
        weight_mem[16'h3618] <= 0;
        weight_mem[16'h3619] <= 0;
        weight_mem[16'h361A] <= 0;
        weight_mem[16'h361B] <= 0;
        weight_mem[16'h361C] <= 0;
        weight_mem[16'h361D] <= 0;
        weight_mem[16'h361E] <= 0;
        weight_mem[16'h361F] <= 0;
        weight_mem[16'h3620] <= 0;
        weight_mem[16'h3621] <= 0;
        weight_mem[16'h3622] <= 0;
        weight_mem[16'h3623] <= 0;
        weight_mem[16'h3624] <= 0;
        weight_mem[16'h3625] <= 0;
        weight_mem[16'h3626] <= 0;
        weight_mem[16'h3627] <= 0;
        weight_mem[16'h3628] <= 0;
        weight_mem[16'h3629] <= 0;
        weight_mem[16'h362A] <= 0;
        weight_mem[16'h362B] <= 0;
        weight_mem[16'h362C] <= 0;
        weight_mem[16'h362D] <= 0;
        weight_mem[16'h362E] <= 0;
        weight_mem[16'h362F] <= 0;
        weight_mem[16'h3630] <= 0;
        weight_mem[16'h3631] <= 0;
        weight_mem[16'h3632] <= 0;
        weight_mem[16'h3633] <= 0;
        weight_mem[16'h3634] <= 0;
        weight_mem[16'h3635] <= 0;
        weight_mem[16'h3636] <= 0;
        weight_mem[16'h3637] <= 0;
        weight_mem[16'h3638] <= 0;
        weight_mem[16'h3639] <= 0;
        weight_mem[16'h363A] <= 0;
        weight_mem[16'h363B] <= 0;
        weight_mem[16'h363C] <= 0;
        weight_mem[16'h363D] <= 0;
        weight_mem[16'h363E] <= 0;
        weight_mem[16'h363F] <= 0;
        weight_mem[16'h3640] <= 0;
        weight_mem[16'h3641] <= 0;
        weight_mem[16'h3642] <= 0;
        weight_mem[16'h3643] <= 0;
        weight_mem[16'h3644] <= 0;
        weight_mem[16'h3645] <= 0;
        weight_mem[16'h3646] <= 0;
        weight_mem[16'h3647] <= 0;
        weight_mem[16'h3648] <= 0;
        weight_mem[16'h3649] <= 0;
        weight_mem[16'h364A] <= 0;
        weight_mem[16'h364B] <= 0;
        weight_mem[16'h364C] <= 0;
        weight_mem[16'h364D] <= 0;
        weight_mem[16'h364E] <= 0;
        weight_mem[16'h364F] <= 0;
        weight_mem[16'h3650] <= 0;
        weight_mem[16'h3651] <= 0;
        weight_mem[16'h3652] <= 0;
        weight_mem[16'h3653] <= 0;
        weight_mem[16'h3654] <= 0;
        weight_mem[16'h3655] <= 0;
        weight_mem[16'h3656] <= 0;
        weight_mem[16'h3657] <= 0;
        weight_mem[16'h3658] <= 0;
        weight_mem[16'h3659] <= 0;
        weight_mem[16'h365A] <= 0;
        weight_mem[16'h365B] <= 0;
        weight_mem[16'h365C] <= 0;
        weight_mem[16'h365D] <= 0;
        weight_mem[16'h365E] <= 0;
        weight_mem[16'h365F] <= 0;
        weight_mem[16'h3660] <= 0;
        weight_mem[16'h3661] <= 0;
        weight_mem[16'h3662] <= 0;
        weight_mem[16'h3663] <= 0;
        weight_mem[16'h3664] <= 0;
        weight_mem[16'h3665] <= 0;
        weight_mem[16'h3666] <= 0;
        weight_mem[16'h3667] <= 0;
        weight_mem[16'h3668] <= 0;
        weight_mem[16'h3669] <= 0;
        weight_mem[16'h366A] <= 0;
        weight_mem[16'h366B] <= 0;
        weight_mem[16'h366C] <= 0;
        weight_mem[16'h366D] <= 0;
        weight_mem[16'h366E] <= 0;
        weight_mem[16'h366F] <= 0;
        weight_mem[16'h3670] <= 0;
        weight_mem[16'h3671] <= 0;
        weight_mem[16'h3672] <= 0;
        weight_mem[16'h3673] <= 0;
        weight_mem[16'h3674] <= 0;
        weight_mem[16'h3675] <= 0;
        weight_mem[16'h3676] <= 0;
        weight_mem[16'h3677] <= 0;
        weight_mem[16'h3678] <= 0;
        weight_mem[16'h3679] <= 0;
        weight_mem[16'h367A] <= 0;
        weight_mem[16'h367B] <= 0;
        weight_mem[16'h367C] <= 0;
        weight_mem[16'h367D] <= 0;
        weight_mem[16'h367E] <= 0;
        weight_mem[16'h367F] <= 0;
        weight_mem[16'h3680] <= 0;
        weight_mem[16'h3681] <= 0;
        weight_mem[16'h3682] <= 0;
        weight_mem[16'h3683] <= 0;
        weight_mem[16'h3684] <= 0;
        weight_mem[16'h3685] <= 0;
        weight_mem[16'h3686] <= 0;
        weight_mem[16'h3687] <= 0;
        weight_mem[16'h3688] <= 0;
        weight_mem[16'h3689] <= 0;
        weight_mem[16'h368A] <= 0;
        weight_mem[16'h368B] <= 0;
        weight_mem[16'h368C] <= 0;
        weight_mem[16'h368D] <= 0;
        weight_mem[16'h368E] <= 0;
        weight_mem[16'h368F] <= 0;
        weight_mem[16'h3690] <= 0;
        weight_mem[16'h3691] <= 0;
        weight_mem[16'h3692] <= 0;
        weight_mem[16'h3693] <= 0;
        weight_mem[16'h3694] <= 0;
        weight_mem[16'h3695] <= 0;
        weight_mem[16'h3696] <= 0;
        weight_mem[16'h3697] <= 0;
        weight_mem[16'h3698] <= 0;
        weight_mem[16'h3699] <= 0;
        weight_mem[16'h369A] <= 0;
        weight_mem[16'h369B] <= 0;
        weight_mem[16'h369C] <= 0;
        weight_mem[16'h369D] <= 0;
        weight_mem[16'h369E] <= 0;
        weight_mem[16'h369F] <= 0;
        weight_mem[16'h36A0] <= 0;
        weight_mem[16'h36A1] <= 0;
        weight_mem[16'h36A2] <= 0;
        weight_mem[16'h36A3] <= 0;
        weight_mem[16'h36A4] <= 0;
        weight_mem[16'h36A5] <= 0;
        weight_mem[16'h36A6] <= 0;
        weight_mem[16'h36A7] <= 0;
        weight_mem[16'h36A8] <= 0;
        weight_mem[16'h36A9] <= 0;
        weight_mem[16'h36AA] <= 0;
        weight_mem[16'h36AB] <= 0;
        weight_mem[16'h36AC] <= 0;
        weight_mem[16'h36AD] <= 0;
        weight_mem[16'h36AE] <= 0;
        weight_mem[16'h36AF] <= 0;
        weight_mem[16'h36B0] <= 0;
        weight_mem[16'h36B1] <= 0;
        weight_mem[16'h36B2] <= 0;
        weight_mem[16'h36B3] <= 0;
        weight_mem[16'h36B4] <= 0;
        weight_mem[16'h36B5] <= 0;
        weight_mem[16'h36B6] <= 0;
        weight_mem[16'h36B7] <= 0;
        weight_mem[16'h36B8] <= 0;
        weight_mem[16'h36B9] <= 0;
        weight_mem[16'h36BA] <= 0;
        weight_mem[16'h36BB] <= 0;
        weight_mem[16'h36BC] <= 0;
        weight_mem[16'h36BD] <= 0;
        weight_mem[16'h36BE] <= 0;
        weight_mem[16'h36BF] <= 0;
        weight_mem[16'h36C0] <= 0;
        weight_mem[16'h36C1] <= 0;
        weight_mem[16'h36C2] <= 0;
        weight_mem[16'h36C3] <= 0;
        weight_mem[16'h36C4] <= 0;
        weight_mem[16'h36C5] <= 0;
        weight_mem[16'h36C6] <= 0;
        weight_mem[16'h36C7] <= 0;
        weight_mem[16'h36C8] <= 0;
        weight_mem[16'h36C9] <= 0;
        weight_mem[16'h36CA] <= 0;
        weight_mem[16'h36CB] <= 0;
        weight_mem[16'h36CC] <= 0;
        weight_mem[16'h36CD] <= 0;
        weight_mem[16'h36CE] <= 0;
        weight_mem[16'h36CF] <= 0;
        weight_mem[16'h36D0] <= 0;
        weight_mem[16'h36D1] <= 0;
        weight_mem[16'h36D2] <= 0;
        weight_mem[16'h36D3] <= 0;
        weight_mem[16'h36D4] <= 0;
        weight_mem[16'h36D5] <= 0;
        weight_mem[16'h36D6] <= 0;
        weight_mem[16'h36D7] <= 0;
        weight_mem[16'h36D8] <= 0;
        weight_mem[16'h36D9] <= 0;
        weight_mem[16'h36DA] <= 0;
        weight_mem[16'h36DB] <= 0;
        weight_mem[16'h36DC] <= 0;
        weight_mem[16'h36DD] <= 0;
        weight_mem[16'h36DE] <= 0;
        weight_mem[16'h36DF] <= 0;
        weight_mem[16'h36E0] <= 0;
        weight_mem[16'h36E1] <= 0;
        weight_mem[16'h36E2] <= 0;
        weight_mem[16'h36E3] <= 0;
        weight_mem[16'h36E4] <= 0;
        weight_mem[16'h36E5] <= 0;
        weight_mem[16'h36E6] <= 0;
        weight_mem[16'h36E7] <= 0;
        weight_mem[16'h36E8] <= 0;
        weight_mem[16'h36E9] <= 0;
        weight_mem[16'h36EA] <= 0;
        weight_mem[16'h36EB] <= 0;
        weight_mem[16'h36EC] <= 0;
        weight_mem[16'h36ED] <= 0;
        weight_mem[16'h36EE] <= 0;
        weight_mem[16'h36EF] <= 0;
        weight_mem[16'h36F0] <= 0;
        weight_mem[16'h36F1] <= 0;
        weight_mem[16'h36F2] <= 0;
        weight_mem[16'h36F3] <= 0;
        weight_mem[16'h36F4] <= 0;
        weight_mem[16'h36F5] <= 0;
        weight_mem[16'h36F6] <= 0;
        weight_mem[16'h36F7] <= 0;
        weight_mem[16'h36F8] <= 0;
        weight_mem[16'h36F9] <= 0;
        weight_mem[16'h36FA] <= 0;
        weight_mem[16'h36FB] <= 0;
        weight_mem[16'h36FC] <= 0;
        weight_mem[16'h36FD] <= 0;
        weight_mem[16'h36FE] <= 0;
        weight_mem[16'h36FF] <= 0;
        weight_mem[16'h3700] <= 0;
        weight_mem[16'h3701] <= 0;
        weight_mem[16'h3702] <= 0;
        weight_mem[16'h3703] <= 0;
        weight_mem[16'h3704] <= 0;
        weight_mem[16'h3705] <= 0;
        weight_mem[16'h3706] <= 0;
        weight_mem[16'h3707] <= 0;
        weight_mem[16'h3708] <= 0;
        weight_mem[16'h3709] <= 0;
        weight_mem[16'h370A] <= 0;
        weight_mem[16'h370B] <= 0;
        weight_mem[16'h370C] <= 0;
        weight_mem[16'h370D] <= 0;
        weight_mem[16'h370E] <= 0;
        weight_mem[16'h370F] <= 0;
        weight_mem[16'h3710] <= 0;
        weight_mem[16'h3711] <= 0;
        weight_mem[16'h3712] <= 0;
        weight_mem[16'h3713] <= 0;
        weight_mem[16'h3714] <= 0;
        weight_mem[16'h3715] <= 0;
        weight_mem[16'h3716] <= 0;
        weight_mem[16'h3717] <= 0;
        weight_mem[16'h3718] <= 0;
        weight_mem[16'h3719] <= 0;
        weight_mem[16'h371A] <= 0;
        weight_mem[16'h371B] <= 0;
        weight_mem[16'h371C] <= 0;
        weight_mem[16'h371D] <= 0;
        weight_mem[16'h371E] <= 0;
        weight_mem[16'h371F] <= 0;
        weight_mem[16'h3720] <= 0;
        weight_mem[16'h3721] <= 0;
        weight_mem[16'h3722] <= 0;
        weight_mem[16'h3723] <= 0;
        weight_mem[16'h3724] <= 0;
        weight_mem[16'h3725] <= 0;
        weight_mem[16'h3726] <= 0;
        weight_mem[16'h3727] <= 0;
        weight_mem[16'h3728] <= 0;
        weight_mem[16'h3729] <= 0;
        weight_mem[16'h372A] <= 0;
        weight_mem[16'h372B] <= 0;
        weight_mem[16'h372C] <= 0;
        weight_mem[16'h372D] <= 0;
        weight_mem[16'h372E] <= 0;
        weight_mem[16'h372F] <= 0;
        weight_mem[16'h3730] <= 0;
        weight_mem[16'h3731] <= 0;
        weight_mem[16'h3732] <= 0;
        weight_mem[16'h3733] <= 0;
        weight_mem[16'h3734] <= 0;
        weight_mem[16'h3735] <= 0;
        weight_mem[16'h3736] <= 0;
        weight_mem[16'h3737] <= 0;
        weight_mem[16'h3738] <= 0;
        weight_mem[16'h3739] <= 0;
        weight_mem[16'h373A] <= 0;
        weight_mem[16'h373B] <= 0;
        weight_mem[16'h373C] <= 0;
        weight_mem[16'h373D] <= 0;
        weight_mem[16'h373E] <= 0;
        weight_mem[16'h373F] <= 0;
        weight_mem[16'h3740] <= 0;
        weight_mem[16'h3741] <= 0;
        weight_mem[16'h3742] <= 0;
        weight_mem[16'h3743] <= 0;
        weight_mem[16'h3744] <= 0;
        weight_mem[16'h3745] <= 0;
        weight_mem[16'h3746] <= 0;
        weight_mem[16'h3747] <= 0;
        weight_mem[16'h3748] <= 0;
        weight_mem[16'h3749] <= 0;
        weight_mem[16'h374A] <= 0;
        weight_mem[16'h374B] <= 0;
        weight_mem[16'h374C] <= 0;
        weight_mem[16'h374D] <= 0;
        weight_mem[16'h374E] <= 0;
        weight_mem[16'h374F] <= 0;
        weight_mem[16'h3750] <= 0;
        weight_mem[16'h3751] <= 0;
        weight_mem[16'h3752] <= 0;
        weight_mem[16'h3753] <= 0;
        weight_mem[16'h3754] <= 0;
        weight_mem[16'h3755] <= 0;
        weight_mem[16'h3756] <= 0;
        weight_mem[16'h3757] <= 0;
        weight_mem[16'h3758] <= 0;
        weight_mem[16'h3759] <= 0;
        weight_mem[16'h375A] <= 0;
        weight_mem[16'h375B] <= 0;
        weight_mem[16'h375C] <= 0;
        weight_mem[16'h375D] <= 0;
        weight_mem[16'h375E] <= 0;
        weight_mem[16'h375F] <= 0;
        weight_mem[16'h3760] <= 0;
        weight_mem[16'h3761] <= 0;
        weight_mem[16'h3762] <= 0;
        weight_mem[16'h3763] <= 0;
        weight_mem[16'h3764] <= 0;
        weight_mem[16'h3765] <= 0;
        weight_mem[16'h3766] <= 0;
        weight_mem[16'h3767] <= 0;
        weight_mem[16'h3768] <= 0;
        weight_mem[16'h3769] <= 0;
        weight_mem[16'h376A] <= 0;
        weight_mem[16'h376B] <= 0;
        weight_mem[16'h376C] <= 0;
        weight_mem[16'h376D] <= 0;
        weight_mem[16'h376E] <= 0;
        weight_mem[16'h376F] <= 0;
        weight_mem[16'h3770] <= 0;
        weight_mem[16'h3771] <= 0;
        weight_mem[16'h3772] <= 0;
        weight_mem[16'h3773] <= 0;
        weight_mem[16'h3774] <= 0;
        weight_mem[16'h3775] <= 0;
        weight_mem[16'h3776] <= 0;
        weight_mem[16'h3777] <= 0;
        weight_mem[16'h3778] <= 0;
        weight_mem[16'h3779] <= 0;
        weight_mem[16'h377A] <= 0;
        weight_mem[16'h377B] <= 0;
        weight_mem[16'h377C] <= 0;
        weight_mem[16'h377D] <= 0;
        weight_mem[16'h377E] <= 0;
        weight_mem[16'h377F] <= 0;
        weight_mem[16'h3780] <= 0;
        weight_mem[16'h3781] <= 0;
        weight_mem[16'h3782] <= 0;
        weight_mem[16'h3783] <= 0;
        weight_mem[16'h3784] <= 0;
        weight_mem[16'h3785] <= 0;
        weight_mem[16'h3786] <= 0;
        weight_mem[16'h3787] <= 0;
        weight_mem[16'h3788] <= 0;
        weight_mem[16'h3789] <= 0;
        weight_mem[16'h378A] <= 0;
        weight_mem[16'h378B] <= 0;
        weight_mem[16'h378C] <= 0;
        weight_mem[16'h378D] <= 0;
        weight_mem[16'h378E] <= 0;
        weight_mem[16'h378F] <= 0;
        weight_mem[16'h3790] <= 0;
        weight_mem[16'h3791] <= 0;
        weight_mem[16'h3792] <= 0;
        weight_mem[16'h3793] <= 0;
        weight_mem[16'h3794] <= 0;
        weight_mem[16'h3795] <= 0;
        weight_mem[16'h3796] <= 0;
        weight_mem[16'h3797] <= 0;
        weight_mem[16'h3798] <= 0;
        weight_mem[16'h3799] <= 0;
        weight_mem[16'h379A] <= 0;
        weight_mem[16'h379B] <= 0;
        weight_mem[16'h379C] <= 0;
        weight_mem[16'h379D] <= 0;
        weight_mem[16'h379E] <= 0;
        weight_mem[16'h379F] <= 0;
        weight_mem[16'h37A0] <= 0;
        weight_mem[16'h37A1] <= 0;
        weight_mem[16'h37A2] <= 0;
        weight_mem[16'h37A3] <= 0;
        weight_mem[16'h37A4] <= 0;
        weight_mem[16'h37A5] <= 0;
        weight_mem[16'h37A6] <= 0;
        weight_mem[16'h37A7] <= 0;
        weight_mem[16'h37A8] <= 0;
        weight_mem[16'h37A9] <= 0;
        weight_mem[16'h37AA] <= 0;
        weight_mem[16'h37AB] <= 0;
        weight_mem[16'h37AC] <= 0;
        weight_mem[16'h37AD] <= 0;
        weight_mem[16'h37AE] <= 0;
        weight_mem[16'h37AF] <= 0;

        // layer 1 neuron 28
        weight_mem[16'h3800] <= 0;
        weight_mem[16'h3801] <= 0;
        weight_mem[16'h3802] <= 0;
        weight_mem[16'h3803] <= 0;
        weight_mem[16'h3804] <= 0;
        weight_mem[16'h3805] <= 0;
        weight_mem[16'h3806] <= 0;
        weight_mem[16'h3807] <= 0;
        weight_mem[16'h3808] <= 0;
        weight_mem[16'h3809] <= 0;
        weight_mem[16'h380A] <= 0;
        weight_mem[16'h380B] <= 0;
        weight_mem[16'h380C] <= 0;
        weight_mem[16'h380D] <= 0;
        weight_mem[16'h380E] <= 0;
        weight_mem[16'h380F] <= 0;
        weight_mem[16'h3810] <= 0;
        weight_mem[16'h3811] <= 0;
        weight_mem[16'h3812] <= 0;
        weight_mem[16'h3813] <= 0;
        weight_mem[16'h3814] <= 0;
        weight_mem[16'h3815] <= 0;
        weight_mem[16'h3816] <= 0;
        weight_mem[16'h3817] <= 0;
        weight_mem[16'h3818] <= 0;
        weight_mem[16'h3819] <= 0;
        weight_mem[16'h381A] <= 0;
        weight_mem[16'h381B] <= 0;
        weight_mem[16'h381C] <= 0;
        weight_mem[16'h381D] <= 0;
        weight_mem[16'h381E] <= 0;
        weight_mem[16'h381F] <= 0;
        weight_mem[16'h3820] <= 0;
        weight_mem[16'h3821] <= 0;
        weight_mem[16'h3822] <= 0;
        weight_mem[16'h3823] <= 0;
        weight_mem[16'h3824] <= 0;
        weight_mem[16'h3825] <= 0;
        weight_mem[16'h3826] <= 0;
        weight_mem[16'h3827] <= 0;
        weight_mem[16'h3828] <= 0;
        weight_mem[16'h3829] <= 0;
        weight_mem[16'h382A] <= 0;
        weight_mem[16'h382B] <= 0;
        weight_mem[16'h382C] <= 0;
        weight_mem[16'h382D] <= 0;
        weight_mem[16'h382E] <= 0;
        weight_mem[16'h382F] <= 0;
        weight_mem[16'h3830] <= 0;
        weight_mem[16'h3831] <= 0;
        weight_mem[16'h3832] <= 0;
        weight_mem[16'h3833] <= 0;
        weight_mem[16'h3834] <= 0;
        weight_mem[16'h3835] <= 0;
        weight_mem[16'h3836] <= 0;
        weight_mem[16'h3837] <= 0;
        weight_mem[16'h3838] <= 0;
        weight_mem[16'h3839] <= 0;
        weight_mem[16'h383A] <= 0;
        weight_mem[16'h383B] <= 0;
        weight_mem[16'h383C] <= 0;
        weight_mem[16'h383D] <= 0;
        weight_mem[16'h383E] <= 0;
        weight_mem[16'h383F] <= 0;
        weight_mem[16'h3840] <= 0;
        weight_mem[16'h3841] <= 0;
        weight_mem[16'h3842] <= 0;
        weight_mem[16'h3843] <= 0;
        weight_mem[16'h3844] <= 0;
        weight_mem[16'h3845] <= 0;
        weight_mem[16'h3846] <= 0;
        weight_mem[16'h3847] <= 0;
        weight_mem[16'h3848] <= 0;
        weight_mem[16'h3849] <= 0;
        weight_mem[16'h384A] <= 0;
        weight_mem[16'h384B] <= 0;
        weight_mem[16'h384C] <= 0;
        weight_mem[16'h384D] <= 0;
        weight_mem[16'h384E] <= 0;
        weight_mem[16'h384F] <= 0;
        weight_mem[16'h3850] <= 0;
        weight_mem[16'h3851] <= 0;
        weight_mem[16'h3852] <= 0;
        weight_mem[16'h3853] <= 0;
        weight_mem[16'h3854] <= 0;
        weight_mem[16'h3855] <= 0;
        weight_mem[16'h3856] <= 0;
        weight_mem[16'h3857] <= 0;
        weight_mem[16'h3858] <= 0;
        weight_mem[16'h3859] <= 0;
        weight_mem[16'h385A] <= 0;
        weight_mem[16'h385B] <= 0;
        weight_mem[16'h385C] <= 0;
        weight_mem[16'h385D] <= 0;
        weight_mem[16'h385E] <= 0;
        weight_mem[16'h385F] <= 0;
        weight_mem[16'h3860] <= 0;
        weight_mem[16'h3861] <= 0;
        weight_mem[16'h3862] <= 0;
        weight_mem[16'h3863] <= 0;
        weight_mem[16'h3864] <= 0;
        weight_mem[16'h3865] <= 0;
        weight_mem[16'h3866] <= 0;
        weight_mem[16'h3867] <= 0;
        weight_mem[16'h3868] <= 0;
        weight_mem[16'h3869] <= 0;
        weight_mem[16'h386A] <= 0;
        weight_mem[16'h386B] <= 0;
        weight_mem[16'h386C] <= 0;
        weight_mem[16'h386D] <= 0;
        weight_mem[16'h386E] <= 0;
        weight_mem[16'h386F] <= 0;
        weight_mem[16'h3870] <= 0;
        weight_mem[16'h3871] <= 0;
        weight_mem[16'h3872] <= 0;
        weight_mem[16'h3873] <= 0;
        weight_mem[16'h3874] <= 0;
        weight_mem[16'h3875] <= 0;
        weight_mem[16'h3876] <= 0;
        weight_mem[16'h3877] <= 0;
        weight_mem[16'h3878] <= 0;
        weight_mem[16'h3879] <= 0;
        weight_mem[16'h387A] <= 0;
        weight_mem[16'h387B] <= 0;
        weight_mem[16'h387C] <= 0;
        weight_mem[16'h387D] <= 0;
        weight_mem[16'h387E] <= 0;
        weight_mem[16'h387F] <= 0;
        weight_mem[16'h3880] <= 0;
        weight_mem[16'h3881] <= 0;
        weight_mem[16'h3882] <= 0;
        weight_mem[16'h3883] <= 0;
        weight_mem[16'h3884] <= 0;
        weight_mem[16'h3885] <= 0;
        weight_mem[16'h3886] <= 0;
        weight_mem[16'h3887] <= 0;
        weight_mem[16'h3888] <= 0;
        weight_mem[16'h3889] <= 0;
        weight_mem[16'h388A] <= 0;
        weight_mem[16'h388B] <= 0;
        weight_mem[16'h388C] <= 0;
        weight_mem[16'h388D] <= 0;
        weight_mem[16'h388E] <= 0;
        weight_mem[16'h388F] <= 0;
        weight_mem[16'h3890] <= 0;
        weight_mem[16'h3891] <= 0;
        weight_mem[16'h3892] <= 0;
        weight_mem[16'h3893] <= 0;
        weight_mem[16'h3894] <= 0;
        weight_mem[16'h3895] <= 0;
        weight_mem[16'h3896] <= 0;
        weight_mem[16'h3897] <= 0;
        weight_mem[16'h3898] <= 0;
        weight_mem[16'h3899] <= 0;
        weight_mem[16'h389A] <= 0;
        weight_mem[16'h389B] <= 0;
        weight_mem[16'h389C] <= 0;
        weight_mem[16'h389D] <= 0;
        weight_mem[16'h389E] <= 0;
        weight_mem[16'h389F] <= 0;
        weight_mem[16'h38A0] <= 0;
        weight_mem[16'h38A1] <= 0;
        weight_mem[16'h38A2] <= 0;
        weight_mem[16'h38A3] <= 0;
        weight_mem[16'h38A4] <= 0;
        weight_mem[16'h38A5] <= 0;
        weight_mem[16'h38A6] <= 0;
        weight_mem[16'h38A7] <= 0;
        weight_mem[16'h38A8] <= 0;
        weight_mem[16'h38A9] <= 0;
        weight_mem[16'h38AA] <= 0;
        weight_mem[16'h38AB] <= 0;
        weight_mem[16'h38AC] <= 0;
        weight_mem[16'h38AD] <= 0;
        weight_mem[16'h38AE] <= 0;
        weight_mem[16'h38AF] <= 0;
        weight_mem[16'h38B0] <= 0;
        weight_mem[16'h38B1] <= 0;
        weight_mem[16'h38B2] <= 0;
        weight_mem[16'h38B3] <= 0;
        weight_mem[16'h38B4] <= 0;
        weight_mem[16'h38B5] <= 0;
        weight_mem[16'h38B6] <= 0;
        weight_mem[16'h38B7] <= 0;
        weight_mem[16'h38B8] <= 0;
        weight_mem[16'h38B9] <= 0;
        weight_mem[16'h38BA] <= 0;
        weight_mem[16'h38BB] <= 0;
        weight_mem[16'h38BC] <= 0;
        weight_mem[16'h38BD] <= 0;
        weight_mem[16'h38BE] <= 0;
        weight_mem[16'h38BF] <= 0;
        weight_mem[16'h38C0] <= 0;
        weight_mem[16'h38C1] <= 0;
        weight_mem[16'h38C2] <= 0;
        weight_mem[16'h38C3] <= 0;
        weight_mem[16'h38C4] <= 0;
        weight_mem[16'h38C5] <= 0;
        weight_mem[16'h38C6] <= 0;
        weight_mem[16'h38C7] <= 0;
        weight_mem[16'h38C8] <= 0;
        weight_mem[16'h38C9] <= 0;
        weight_mem[16'h38CA] <= 0;
        weight_mem[16'h38CB] <= 0;
        weight_mem[16'h38CC] <= 0;
        weight_mem[16'h38CD] <= 0;
        weight_mem[16'h38CE] <= 0;
        weight_mem[16'h38CF] <= 0;
        weight_mem[16'h38D0] <= 0;
        weight_mem[16'h38D1] <= 0;
        weight_mem[16'h38D2] <= 0;
        weight_mem[16'h38D3] <= 0;
        weight_mem[16'h38D4] <= 0;
        weight_mem[16'h38D5] <= 0;
        weight_mem[16'h38D6] <= 0;
        weight_mem[16'h38D7] <= 0;
        weight_mem[16'h38D8] <= 0;
        weight_mem[16'h38D9] <= 0;
        weight_mem[16'h38DA] <= 0;
        weight_mem[16'h38DB] <= 0;
        weight_mem[16'h38DC] <= 0;
        weight_mem[16'h38DD] <= 0;
        weight_mem[16'h38DE] <= 0;
        weight_mem[16'h38DF] <= 0;
        weight_mem[16'h38E0] <= 0;
        weight_mem[16'h38E1] <= 0;
        weight_mem[16'h38E2] <= 0;
        weight_mem[16'h38E3] <= 0;
        weight_mem[16'h38E4] <= 0;
        weight_mem[16'h38E5] <= 0;
        weight_mem[16'h38E6] <= 0;
        weight_mem[16'h38E7] <= 0;
        weight_mem[16'h38E8] <= 0;
        weight_mem[16'h38E9] <= 0;
        weight_mem[16'h38EA] <= 0;
        weight_mem[16'h38EB] <= 0;
        weight_mem[16'h38EC] <= 0;
        weight_mem[16'h38ED] <= 0;
        weight_mem[16'h38EE] <= 0;
        weight_mem[16'h38EF] <= 0;
        weight_mem[16'h38F0] <= 0;
        weight_mem[16'h38F1] <= 0;
        weight_mem[16'h38F2] <= 0;
        weight_mem[16'h38F3] <= 0;
        weight_mem[16'h38F4] <= 0;
        weight_mem[16'h38F5] <= 0;
        weight_mem[16'h38F6] <= 0;
        weight_mem[16'h38F7] <= 0;
        weight_mem[16'h38F8] <= 0;
        weight_mem[16'h38F9] <= 0;
        weight_mem[16'h38FA] <= 0;
        weight_mem[16'h38FB] <= 0;
        weight_mem[16'h38FC] <= 0;
        weight_mem[16'h38FD] <= 0;
        weight_mem[16'h38FE] <= 0;
        weight_mem[16'h38FF] <= 0;
        weight_mem[16'h3900] <= 0;
        weight_mem[16'h3901] <= 0;
        weight_mem[16'h3902] <= 0;
        weight_mem[16'h3903] <= 0;
        weight_mem[16'h3904] <= 0;
        weight_mem[16'h3905] <= 0;
        weight_mem[16'h3906] <= 0;
        weight_mem[16'h3907] <= 0;
        weight_mem[16'h3908] <= 0;
        weight_mem[16'h3909] <= 0;
        weight_mem[16'h390A] <= 0;
        weight_mem[16'h390B] <= 0;
        weight_mem[16'h390C] <= 0;
        weight_mem[16'h390D] <= 0;
        weight_mem[16'h390E] <= 0;
        weight_mem[16'h390F] <= 0;
        weight_mem[16'h3910] <= 0;
        weight_mem[16'h3911] <= 0;
        weight_mem[16'h3912] <= 0;
        weight_mem[16'h3913] <= 0;
        weight_mem[16'h3914] <= 0;
        weight_mem[16'h3915] <= 0;
        weight_mem[16'h3916] <= 0;
        weight_mem[16'h3917] <= 0;
        weight_mem[16'h3918] <= 0;
        weight_mem[16'h3919] <= 0;
        weight_mem[16'h391A] <= 0;
        weight_mem[16'h391B] <= 0;
        weight_mem[16'h391C] <= 0;
        weight_mem[16'h391D] <= 0;
        weight_mem[16'h391E] <= 0;
        weight_mem[16'h391F] <= 0;
        weight_mem[16'h3920] <= 0;
        weight_mem[16'h3921] <= 0;
        weight_mem[16'h3922] <= 0;
        weight_mem[16'h3923] <= 0;
        weight_mem[16'h3924] <= 0;
        weight_mem[16'h3925] <= 0;
        weight_mem[16'h3926] <= 0;
        weight_mem[16'h3927] <= 0;
        weight_mem[16'h3928] <= 0;
        weight_mem[16'h3929] <= 0;
        weight_mem[16'h392A] <= 0;
        weight_mem[16'h392B] <= 0;
        weight_mem[16'h392C] <= 0;
        weight_mem[16'h392D] <= 0;
        weight_mem[16'h392E] <= 0;
        weight_mem[16'h392F] <= 0;
        weight_mem[16'h3930] <= 0;
        weight_mem[16'h3931] <= 0;
        weight_mem[16'h3932] <= 0;
        weight_mem[16'h3933] <= 0;
        weight_mem[16'h3934] <= 0;
        weight_mem[16'h3935] <= 0;
        weight_mem[16'h3936] <= 0;
        weight_mem[16'h3937] <= 0;
        weight_mem[16'h3938] <= 0;
        weight_mem[16'h3939] <= 0;
        weight_mem[16'h393A] <= 0;
        weight_mem[16'h393B] <= 0;
        weight_mem[16'h393C] <= 0;
        weight_mem[16'h393D] <= 0;
        weight_mem[16'h393E] <= 0;
        weight_mem[16'h393F] <= 0;
        weight_mem[16'h3940] <= 0;
        weight_mem[16'h3941] <= 0;
        weight_mem[16'h3942] <= 0;
        weight_mem[16'h3943] <= 0;
        weight_mem[16'h3944] <= 0;
        weight_mem[16'h3945] <= 0;
        weight_mem[16'h3946] <= 0;
        weight_mem[16'h3947] <= 0;
        weight_mem[16'h3948] <= 0;
        weight_mem[16'h3949] <= 0;
        weight_mem[16'h394A] <= 0;
        weight_mem[16'h394B] <= 0;
        weight_mem[16'h394C] <= 0;
        weight_mem[16'h394D] <= 0;
        weight_mem[16'h394E] <= 0;
        weight_mem[16'h394F] <= 0;
        weight_mem[16'h3950] <= 0;
        weight_mem[16'h3951] <= 0;
        weight_mem[16'h3952] <= 0;
        weight_mem[16'h3953] <= 0;
        weight_mem[16'h3954] <= 0;
        weight_mem[16'h3955] <= 0;
        weight_mem[16'h3956] <= 0;
        weight_mem[16'h3957] <= 0;
        weight_mem[16'h3958] <= 0;
        weight_mem[16'h3959] <= 0;
        weight_mem[16'h395A] <= 0;
        weight_mem[16'h395B] <= 0;
        weight_mem[16'h395C] <= 0;
        weight_mem[16'h395D] <= 0;
        weight_mem[16'h395E] <= 0;
        weight_mem[16'h395F] <= 0;
        weight_mem[16'h3960] <= 0;
        weight_mem[16'h3961] <= 0;
        weight_mem[16'h3962] <= 0;
        weight_mem[16'h3963] <= 0;
        weight_mem[16'h3964] <= 0;
        weight_mem[16'h3965] <= 0;
        weight_mem[16'h3966] <= 0;
        weight_mem[16'h3967] <= 0;
        weight_mem[16'h3968] <= 0;
        weight_mem[16'h3969] <= 0;
        weight_mem[16'h396A] <= 0;
        weight_mem[16'h396B] <= 0;
        weight_mem[16'h396C] <= 0;
        weight_mem[16'h396D] <= 0;
        weight_mem[16'h396E] <= 0;
        weight_mem[16'h396F] <= 0;
        weight_mem[16'h3970] <= 0;
        weight_mem[16'h3971] <= 0;
        weight_mem[16'h3972] <= 0;
        weight_mem[16'h3973] <= 0;
        weight_mem[16'h3974] <= 0;
        weight_mem[16'h3975] <= 0;
        weight_mem[16'h3976] <= 0;
        weight_mem[16'h3977] <= 0;
        weight_mem[16'h3978] <= 0;
        weight_mem[16'h3979] <= 0;
        weight_mem[16'h397A] <= 0;
        weight_mem[16'h397B] <= 0;
        weight_mem[16'h397C] <= 0;
        weight_mem[16'h397D] <= 0;
        weight_mem[16'h397E] <= 0;
        weight_mem[16'h397F] <= 0;
        weight_mem[16'h3980] <= 0;
        weight_mem[16'h3981] <= 0;
        weight_mem[16'h3982] <= 0;
        weight_mem[16'h3983] <= 0;
        weight_mem[16'h3984] <= 0;
        weight_mem[16'h3985] <= 0;
        weight_mem[16'h3986] <= 0;
        weight_mem[16'h3987] <= 0;
        weight_mem[16'h3988] <= 0;
        weight_mem[16'h3989] <= 0;
        weight_mem[16'h398A] <= 0;
        weight_mem[16'h398B] <= 0;
        weight_mem[16'h398C] <= 0;
        weight_mem[16'h398D] <= 0;
        weight_mem[16'h398E] <= 0;
        weight_mem[16'h398F] <= 0;
        weight_mem[16'h3990] <= 0;
        weight_mem[16'h3991] <= 0;
        weight_mem[16'h3992] <= 0;
        weight_mem[16'h3993] <= 0;
        weight_mem[16'h3994] <= 0;
        weight_mem[16'h3995] <= 0;
        weight_mem[16'h3996] <= 0;
        weight_mem[16'h3997] <= 0;
        weight_mem[16'h3998] <= 0;
        weight_mem[16'h3999] <= 0;
        weight_mem[16'h399A] <= 0;
        weight_mem[16'h399B] <= 0;
        weight_mem[16'h399C] <= 0;
        weight_mem[16'h399D] <= 0;
        weight_mem[16'h399E] <= 0;
        weight_mem[16'h399F] <= 0;
        weight_mem[16'h39A0] <= 0;
        weight_mem[16'h39A1] <= 0;
        weight_mem[16'h39A2] <= 0;
        weight_mem[16'h39A3] <= 0;
        weight_mem[16'h39A4] <= 0;
        weight_mem[16'h39A5] <= 0;
        weight_mem[16'h39A6] <= 0;
        weight_mem[16'h39A7] <= 0;
        weight_mem[16'h39A8] <= 0;
        weight_mem[16'h39A9] <= 0;
        weight_mem[16'h39AA] <= 0;
        weight_mem[16'h39AB] <= 0;
        weight_mem[16'h39AC] <= 0;
        weight_mem[16'h39AD] <= 0;
        weight_mem[16'h39AE] <= 0;
        weight_mem[16'h39AF] <= 0;

        // layer 1 neuron 29
        weight_mem[16'h3A00] <= 0;
        weight_mem[16'h3A01] <= 0;
        weight_mem[16'h3A02] <= 0;
        weight_mem[16'h3A03] <= 0;
        weight_mem[16'h3A04] <= 0;
        weight_mem[16'h3A05] <= 0;
        weight_mem[16'h3A06] <= 0;
        weight_mem[16'h3A07] <= 0;
        weight_mem[16'h3A08] <= 0;
        weight_mem[16'h3A09] <= 0;
        weight_mem[16'h3A0A] <= 0;
        weight_mem[16'h3A0B] <= 0;
        weight_mem[16'h3A0C] <= 0;
        weight_mem[16'h3A0D] <= 0;
        weight_mem[16'h3A0E] <= 0;
        weight_mem[16'h3A0F] <= 0;
        weight_mem[16'h3A10] <= 0;
        weight_mem[16'h3A11] <= 0;
        weight_mem[16'h3A12] <= 0;
        weight_mem[16'h3A13] <= 0;
        weight_mem[16'h3A14] <= 0;
        weight_mem[16'h3A15] <= 0;
        weight_mem[16'h3A16] <= 0;
        weight_mem[16'h3A17] <= 0;
        weight_mem[16'h3A18] <= 0;
        weight_mem[16'h3A19] <= 0;
        weight_mem[16'h3A1A] <= 0;
        weight_mem[16'h3A1B] <= 0;
        weight_mem[16'h3A1C] <= 0;
        weight_mem[16'h3A1D] <= 0;
        weight_mem[16'h3A1E] <= 0;
        weight_mem[16'h3A1F] <= 0;
        weight_mem[16'h3A20] <= 0;
        weight_mem[16'h3A21] <= 0;
        weight_mem[16'h3A22] <= 0;
        weight_mem[16'h3A23] <= 0;
        weight_mem[16'h3A24] <= 0;
        weight_mem[16'h3A25] <= 0;
        weight_mem[16'h3A26] <= 0;
        weight_mem[16'h3A27] <= 0;
        weight_mem[16'h3A28] <= 0;
        weight_mem[16'h3A29] <= 0;
        weight_mem[16'h3A2A] <= 0;
        weight_mem[16'h3A2B] <= 0;
        weight_mem[16'h3A2C] <= 0;
        weight_mem[16'h3A2D] <= 0;
        weight_mem[16'h3A2E] <= 0;
        weight_mem[16'h3A2F] <= 0;
        weight_mem[16'h3A30] <= 0;
        weight_mem[16'h3A31] <= 0;
        weight_mem[16'h3A32] <= 0;
        weight_mem[16'h3A33] <= 0;
        weight_mem[16'h3A34] <= 0;
        weight_mem[16'h3A35] <= 0;
        weight_mem[16'h3A36] <= 0;
        weight_mem[16'h3A37] <= 0;
        weight_mem[16'h3A38] <= 0;
        weight_mem[16'h3A39] <= 0;
        weight_mem[16'h3A3A] <= 0;
        weight_mem[16'h3A3B] <= 0;
        weight_mem[16'h3A3C] <= 0;
        weight_mem[16'h3A3D] <= 0;
        weight_mem[16'h3A3E] <= 0;
        weight_mem[16'h3A3F] <= 0;
        weight_mem[16'h3A40] <= 0;
        weight_mem[16'h3A41] <= 0;
        weight_mem[16'h3A42] <= 0;
        weight_mem[16'h3A43] <= 0;
        weight_mem[16'h3A44] <= 0;
        weight_mem[16'h3A45] <= 0;
        weight_mem[16'h3A46] <= 0;
        weight_mem[16'h3A47] <= 0;
        weight_mem[16'h3A48] <= 0;
        weight_mem[16'h3A49] <= 0;
        weight_mem[16'h3A4A] <= 0;
        weight_mem[16'h3A4B] <= 0;
        weight_mem[16'h3A4C] <= 0;
        weight_mem[16'h3A4D] <= 0;
        weight_mem[16'h3A4E] <= 0;
        weight_mem[16'h3A4F] <= 0;
        weight_mem[16'h3A50] <= 0;
        weight_mem[16'h3A51] <= 0;
        weight_mem[16'h3A52] <= 0;
        weight_mem[16'h3A53] <= 0;
        weight_mem[16'h3A54] <= 0;
        weight_mem[16'h3A55] <= 0;
        weight_mem[16'h3A56] <= 0;
        weight_mem[16'h3A57] <= 0;
        weight_mem[16'h3A58] <= 0;
        weight_mem[16'h3A59] <= 0;
        weight_mem[16'h3A5A] <= 0;
        weight_mem[16'h3A5B] <= 0;
        weight_mem[16'h3A5C] <= 0;
        weight_mem[16'h3A5D] <= 0;
        weight_mem[16'h3A5E] <= 0;
        weight_mem[16'h3A5F] <= 0;
        weight_mem[16'h3A60] <= 0;
        weight_mem[16'h3A61] <= 0;
        weight_mem[16'h3A62] <= 0;
        weight_mem[16'h3A63] <= 0;
        weight_mem[16'h3A64] <= 0;
        weight_mem[16'h3A65] <= 0;
        weight_mem[16'h3A66] <= 0;
        weight_mem[16'h3A67] <= 0;
        weight_mem[16'h3A68] <= 0;
        weight_mem[16'h3A69] <= 0;
        weight_mem[16'h3A6A] <= 0;
        weight_mem[16'h3A6B] <= 0;
        weight_mem[16'h3A6C] <= 0;
        weight_mem[16'h3A6D] <= 0;
        weight_mem[16'h3A6E] <= 0;
        weight_mem[16'h3A6F] <= 0;
        weight_mem[16'h3A70] <= 0;
        weight_mem[16'h3A71] <= 0;
        weight_mem[16'h3A72] <= 0;
        weight_mem[16'h3A73] <= 0;
        weight_mem[16'h3A74] <= 0;
        weight_mem[16'h3A75] <= 0;
        weight_mem[16'h3A76] <= 0;
        weight_mem[16'h3A77] <= 0;
        weight_mem[16'h3A78] <= 0;
        weight_mem[16'h3A79] <= 0;
        weight_mem[16'h3A7A] <= 0;
        weight_mem[16'h3A7B] <= 0;
        weight_mem[16'h3A7C] <= 0;
        weight_mem[16'h3A7D] <= 0;
        weight_mem[16'h3A7E] <= 0;
        weight_mem[16'h3A7F] <= 0;
        weight_mem[16'h3A80] <= 0;
        weight_mem[16'h3A81] <= 0;
        weight_mem[16'h3A82] <= 0;
        weight_mem[16'h3A83] <= 0;
        weight_mem[16'h3A84] <= 0;
        weight_mem[16'h3A85] <= 0;
        weight_mem[16'h3A86] <= 0;
        weight_mem[16'h3A87] <= 0;
        weight_mem[16'h3A88] <= 0;
        weight_mem[16'h3A89] <= 0;
        weight_mem[16'h3A8A] <= 0;
        weight_mem[16'h3A8B] <= 0;
        weight_mem[16'h3A8C] <= 0;
        weight_mem[16'h3A8D] <= 0;
        weight_mem[16'h3A8E] <= 0;
        weight_mem[16'h3A8F] <= 0;
        weight_mem[16'h3A90] <= 0;
        weight_mem[16'h3A91] <= 0;
        weight_mem[16'h3A92] <= 0;
        weight_mem[16'h3A93] <= 0;
        weight_mem[16'h3A94] <= 0;
        weight_mem[16'h3A95] <= 0;
        weight_mem[16'h3A96] <= 0;
        weight_mem[16'h3A97] <= 0;
        weight_mem[16'h3A98] <= 0;
        weight_mem[16'h3A99] <= 0;
        weight_mem[16'h3A9A] <= 0;
        weight_mem[16'h3A9B] <= 0;
        weight_mem[16'h3A9C] <= 0;
        weight_mem[16'h3A9D] <= 0;
        weight_mem[16'h3A9E] <= 0;
        weight_mem[16'h3A9F] <= 0;
        weight_mem[16'h3AA0] <= 0;
        weight_mem[16'h3AA1] <= 0;
        weight_mem[16'h3AA2] <= 0;
        weight_mem[16'h3AA3] <= 0;
        weight_mem[16'h3AA4] <= 0;
        weight_mem[16'h3AA5] <= 0;
        weight_mem[16'h3AA6] <= 0;
        weight_mem[16'h3AA7] <= 0;
        weight_mem[16'h3AA8] <= 0;
        weight_mem[16'h3AA9] <= 0;
        weight_mem[16'h3AAA] <= 0;
        weight_mem[16'h3AAB] <= 0;
        weight_mem[16'h3AAC] <= 0;
        weight_mem[16'h3AAD] <= 0;
        weight_mem[16'h3AAE] <= 0;
        weight_mem[16'h3AAF] <= 0;
        weight_mem[16'h3AB0] <= 0;
        weight_mem[16'h3AB1] <= 0;
        weight_mem[16'h3AB2] <= 0;
        weight_mem[16'h3AB3] <= 0;
        weight_mem[16'h3AB4] <= 0;
        weight_mem[16'h3AB5] <= 0;
        weight_mem[16'h3AB6] <= 0;
        weight_mem[16'h3AB7] <= 0;
        weight_mem[16'h3AB8] <= 0;
        weight_mem[16'h3AB9] <= 0;
        weight_mem[16'h3ABA] <= 0;
        weight_mem[16'h3ABB] <= 0;
        weight_mem[16'h3ABC] <= 0;
        weight_mem[16'h3ABD] <= 0;
        weight_mem[16'h3ABE] <= 0;
        weight_mem[16'h3ABF] <= 0;
        weight_mem[16'h3AC0] <= 0;
        weight_mem[16'h3AC1] <= 0;
        weight_mem[16'h3AC2] <= 0;
        weight_mem[16'h3AC3] <= 0;
        weight_mem[16'h3AC4] <= 0;
        weight_mem[16'h3AC5] <= 0;
        weight_mem[16'h3AC6] <= 0;
        weight_mem[16'h3AC7] <= 0;
        weight_mem[16'h3AC8] <= 0;
        weight_mem[16'h3AC9] <= 0;
        weight_mem[16'h3ACA] <= 0;
        weight_mem[16'h3ACB] <= 0;
        weight_mem[16'h3ACC] <= 0;
        weight_mem[16'h3ACD] <= 0;
        weight_mem[16'h3ACE] <= 0;
        weight_mem[16'h3ACF] <= 0;
        weight_mem[16'h3AD0] <= 0;
        weight_mem[16'h3AD1] <= 0;
        weight_mem[16'h3AD2] <= 0;
        weight_mem[16'h3AD3] <= 0;
        weight_mem[16'h3AD4] <= 0;
        weight_mem[16'h3AD5] <= 0;
        weight_mem[16'h3AD6] <= 0;
        weight_mem[16'h3AD7] <= 0;
        weight_mem[16'h3AD8] <= 0;
        weight_mem[16'h3AD9] <= 0;
        weight_mem[16'h3ADA] <= 0;
        weight_mem[16'h3ADB] <= 0;
        weight_mem[16'h3ADC] <= 0;
        weight_mem[16'h3ADD] <= 0;
        weight_mem[16'h3ADE] <= 0;
        weight_mem[16'h3ADF] <= 0;
        weight_mem[16'h3AE0] <= 0;
        weight_mem[16'h3AE1] <= 0;
        weight_mem[16'h3AE2] <= 0;
        weight_mem[16'h3AE3] <= 0;
        weight_mem[16'h3AE4] <= 0;
        weight_mem[16'h3AE5] <= 0;
        weight_mem[16'h3AE6] <= 0;
        weight_mem[16'h3AE7] <= 0;
        weight_mem[16'h3AE8] <= 0;
        weight_mem[16'h3AE9] <= 0;
        weight_mem[16'h3AEA] <= 0;
        weight_mem[16'h3AEB] <= 0;
        weight_mem[16'h3AEC] <= 0;
        weight_mem[16'h3AED] <= 0;
        weight_mem[16'h3AEE] <= 0;
        weight_mem[16'h3AEF] <= 0;
        weight_mem[16'h3AF0] <= 0;
        weight_mem[16'h3AF1] <= 0;
        weight_mem[16'h3AF2] <= 0;
        weight_mem[16'h3AF3] <= 0;
        weight_mem[16'h3AF4] <= 0;
        weight_mem[16'h3AF5] <= 0;
        weight_mem[16'h3AF6] <= 0;
        weight_mem[16'h3AF7] <= 0;
        weight_mem[16'h3AF8] <= 0;
        weight_mem[16'h3AF9] <= 0;
        weight_mem[16'h3AFA] <= 0;
        weight_mem[16'h3AFB] <= 0;
        weight_mem[16'h3AFC] <= 0;
        weight_mem[16'h3AFD] <= 0;
        weight_mem[16'h3AFE] <= 0;
        weight_mem[16'h3AFF] <= 0;
        weight_mem[16'h3B00] <= 0;
        weight_mem[16'h3B01] <= 0;
        weight_mem[16'h3B02] <= 0;
        weight_mem[16'h3B03] <= 0;
        weight_mem[16'h3B04] <= 0;
        weight_mem[16'h3B05] <= 0;
        weight_mem[16'h3B06] <= 0;
        weight_mem[16'h3B07] <= 0;
        weight_mem[16'h3B08] <= 0;
        weight_mem[16'h3B09] <= 0;
        weight_mem[16'h3B0A] <= 0;
        weight_mem[16'h3B0B] <= 0;
        weight_mem[16'h3B0C] <= 0;
        weight_mem[16'h3B0D] <= 0;
        weight_mem[16'h3B0E] <= 0;
        weight_mem[16'h3B0F] <= 0;
        weight_mem[16'h3B10] <= 0;
        weight_mem[16'h3B11] <= 0;
        weight_mem[16'h3B12] <= 0;
        weight_mem[16'h3B13] <= 0;
        weight_mem[16'h3B14] <= 0;
        weight_mem[16'h3B15] <= 0;
        weight_mem[16'h3B16] <= 0;
        weight_mem[16'h3B17] <= 0;
        weight_mem[16'h3B18] <= 0;
        weight_mem[16'h3B19] <= 0;
        weight_mem[16'h3B1A] <= 0;
        weight_mem[16'h3B1B] <= 0;
        weight_mem[16'h3B1C] <= 0;
        weight_mem[16'h3B1D] <= 0;
        weight_mem[16'h3B1E] <= 0;
        weight_mem[16'h3B1F] <= 0;
        weight_mem[16'h3B20] <= 0;
        weight_mem[16'h3B21] <= 0;
        weight_mem[16'h3B22] <= 0;
        weight_mem[16'h3B23] <= 0;
        weight_mem[16'h3B24] <= 0;
        weight_mem[16'h3B25] <= 0;
        weight_mem[16'h3B26] <= 0;
        weight_mem[16'h3B27] <= 0;
        weight_mem[16'h3B28] <= 0;
        weight_mem[16'h3B29] <= 0;
        weight_mem[16'h3B2A] <= 0;
        weight_mem[16'h3B2B] <= 0;
        weight_mem[16'h3B2C] <= 0;
        weight_mem[16'h3B2D] <= 0;
        weight_mem[16'h3B2E] <= 0;
        weight_mem[16'h3B2F] <= 0;
        weight_mem[16'h3B30] <= 0;
        weight_mem[16'h3B31] <= 0;
        weight_mem[16'h3B32] <= 0;
        weight_mem[16'h3B33] <= 0;
        weight_mem[16'h3B34] <= 0;
        weight_mem[16'h3B35] <= 0;
        weight_mem[16'h3B36] <= 0;
        weight_mem[16'h3B37] <= 0;
        weight_mem[16'h3B38] <= 0;
        weight_mem[16'h3B39] <= 0;
        weight_mem[16'h3B3A] <= 0;
        weight_mem[16'h3B3B] <= 0;
        weight_mem[16'h3B3C] <= 0;
        weight_mem[16'h3B3D] <= 0;
        weight_mem[16'h3B3E] <= 0;
        weight_mem[16'h3B3F] <= 0;
        weight_mem[16'h3B40] <= 0;
        weight_mem[16'h3B41] <= 0;
        weight_mem[16'h3B42] <= 0;
        weight_mem[16'h3B43] <= 0;
        weight_mem[16'h3B44] <= 0;
        weight_mem[16'h3B45] <= 0;
        weight_mem[16'h3B46] <= 0;
        weight_mem[16'h3B47] <= 0;
        weight_mem[16'h3B48] <= 0;
        weight_mem[16'h3B49] <= 0;
        weight_mem[16'h3B4A] <= 0;
        weight_mem[16'h3B4B] <= 0;
        weight_mem[16'h3B4C] <= 0;
        weight_mem[16'h3B4D] <= 0;
        weight_mem[16'h3B4E] <= 0;
        weight_mem[16'h3B4F] <= 0;
        weight_mem[16'h3B50] <= 0;
        weight_mem[16'h3B51] <= 0;
        weight_mem[16'h3B52] <= 0;
        weight_mem[16'h3B53] <= 0;
        weight_mem[16'h3B54] <= 0;
        weight_mem[16'h3B55] <= 0;
        weight_mem[16'h3B56] <= 0;
        weight_mem[16'h3B57] <= 0;
        weight_mem[16'h3B58] <= 0;
        weight_mem[16'h3B59] <= 0;
        weight_mem[16'h3B5A] <= 0;
        weight_mem[16'h3B5B] <= 0;
        weight_mem[16'h3B5C] <= 0;
        weight_mem[16'h3B5D] <= 0;
        weight_mem[16'h3B5E] <= 0;
        weight_mem[16'h3B5F] <= 0;
        weight_mem[16'h3B60] <= 0;
        weight_mem[16'h3B61] <= 0;
        weight_mem[16'h3B62] <= 0;
        weight_mem[16'h3B63] <= 0;
        weight_mem[16'h3B64] <= 0;
        weight_mem[16'h3B65] <= 0;
        weight_mem[16'h3B66] <= 0;
        weight_mem[16'h3B67] <= 0;
        weight_mem[16'h3B68] <= 0;
        weight_mem[16'h3B69] <= 0;
        weight_mem[16'h3B6A] <= 0;
        weight_mem[16'h3B6B] <= 0;
        weight_mem[16'h3B6C] <= 0;
        weight_mem[16'h3B6D] <= 0;
        weight_mem[16'h3B6E] <= 0;
        weight_mem[16'h3B6F] <= 0;
        weight_mem[16'h3B70] <= 0;
        weight_mem[16'h3B71] <= 0;
        weight_mem[16'h3B72] <= 0;
        weight_mem[16'h3B73] <= 0;
        weight_mem[16'h3B74] <= 0;
        weight_mem[16'h3B75] <= 0;
        weight_mem[16'h3B76] <= 0;
        weight_mem[16'h3B77] <= 0;
        weight_mem[16'h3B78] <= 0;
        weight_mem[16'h3B79] <= 0;
        weight_mem[16'h3B7A] <= 0;
        weight_mem[16'h3B7B] <= 0;
        weight_mem[16'h3B7C] <= 0;
        weight_mem[16'h3B7D] <= 0;
        weight_mem[16'h3B7E] <= 0;
        weight_mem[16'h3B7F] <= 0;
        weight_mem[16'h3B80] <= 0;
        weight_mem[16'h3B81] <= 0;
        weight_mem[16'h3B82] <= 0;
        weight_mem[16'h3B83] <= 0;
        weight_mem[16'h3B84] <= 0;
        weight_mem[16'h3B85] <= 0;
        weight_mem[16'h3B86] <= 0;
        weight_mem[16'h3B87] <= 0;
        weight_mem[16'h3B88] <= 0;
        weight_mem[16'h3B89] <= 0;
        weight_mem[16'h3B8A] <= 0;
        weight_mem[16'h3B8B] <= 0;
        weight_mem[16'h3B8C] <= 0;
        weight_mem[16'h3B8D] <= 0;
        weight_mem[16'h3B8E] <= 0;
        weight_mem[16'h3B8F] <= 0;
        weight_mem[16'h3B90] <= 0;
        weight_mem[16'h3B91] <= 0;
        weight_mem[16'h3B92] <= 0;
        weight_mem[16'h3B93] <= 0;
        weight_mem[16'h3B94] <= 0;
        weight_mem[16'h3B95] <= 0;
        weight_mem[16'h3B96] <= 0;
        weight_mem[16'h3B97] <= 0;
        weight_mem[16'h3B98] <= 0;
        weight_mem[16'h3B99] <= 0;
        weight_mem[16'h3B9A] <= 0;
        weight_mem[16'h3B9B] <= 0;
        weight_mem[16'h3B9C] <= 0;
        weight_mem[16'h3B9D] <= 0;
        weight_mem[16'h3B9E] <= 0;
        weight_mem[16'h3B9F] <= 0;
        weight_mem[16'h3BA0] <= 0;
        weight_mem[16'h3BA1] <= 0;
        weight_mem[16'h3BA2] <= 0;
        weight_mem[16'h3BA3] <= 0;
        weight_mem[16'h3BA4] <= 0;
        weight_mem[16'h3BA5] <= 0;
        weight_mem[16'h3BA6] <= 0;
        weight_mem[16'h3BA7] <= 0;
        weight_mem[16'h3BA8] <= 0;
        weight_mem[16'h3BA9] <= 0;
        weight_mem[16'h3BAA] <= 0;
        weight_mem[16'h3BAB] <= 0;
        weight_mem[16'h3BAC] <= 0;
        weight_mem[16'h3BAD] <= 0;
        weight_mem[16'h3BAE] <= 0;
        weight_mem[16'h3BAF] <= 0;

        // layer 2 neuron 0
        weight_mem[16'h4000] <= 1;
        weight_mem[16'h4001] <= 0;
        weight_mem[16'h4002] <= 0;
        weight_mem[16'h4003] <= 0;
        weight_mem[16'h4004] <= 0;
        weight_mem[16'h4005] <= 0;
        weight_mem[16'h4006] <= 0;
        weight_mem[16'h4007] <= 0;
        weight_mem[16'h4008] <= 0;
        weight_mem[16'h4009] <= 0;
        weight_mem[16'h400A] <= 0;
        weight_mem[16'h400B] <= 0;
        weight_mem[16'h400C] <= 0;
        weight_mem[16'h400D] <= 0;
        weight_mem[16'h400E] <= 0;
        weight_mem[16'h400F] <= 0;
        weight_mem[16'h4010] <= 0;
        weight_mem[16'h4011] <= 0;
        weight_mem[16'h4012] <= 0;
        weight_mem[16'h4013] <= 0;
        weight_mem[16'h4014] <= 0;
        weight_mem[16'h4015] <= 0;
        weight_mem[16'h4016] <= 0;
        weight_mem[16'h4017] <= 0;
        weight_mem[16'h4018] <= 0;
        weight_mem[16'h4019] <= 0;
        weight_mem[16'h401A] <= 0;
        weight_mem[16'h401B] <= 0;
        weight_mem[16'h401C] <= 0;
        weight_mem[16'h401D] <= 0;

        // layer 2 neuron 1
        weight_mem[16'h4200] <= 0;
        weight_mem[16'h4201] <= 0;
        weight_mem[16'h4202] <= 0;
        weight_mem[16'h4203] <= 0;
        weight_mem[16'h4204] <= 0;
        weight_mem[16'h4205] <= 0;
        weight_mem[16'h4206] <= 0;
        weight_mem[16'h4207] <= 0;
        weight_mem[16'h4208] <= 0;
        weight_mem[16'h4209] <= 0;
        weight_mem[16'h420A] <= 0;
        weight_mem[16'h420B] <= 0;
        weight_mem[16'h420C] <= 0;
        weight_mem[16'h420D] <= 0;
        weight_mem[16'h420E] <= 0;
        weight_mem[16'h420F] <= 0;
        weight_mem[16'h4210] <= 0;
        weight_mem[16'h4211] <= 0;
        weight_mem[16'h4212] <= 0;
        weight_mem[16'h4213] <= 0;
        weight_mem[16'h4214] <= 0;
        weight_mem[16'h4215] <= 0;
        weight_mem[16'h4216] <= 0;
        weight_mem[16'h4217] <= 0;
        weight_mem[16'h4218] <= 0;
        weight_mem[16'h4219] <= 0;
        weight_mem[16'h421A] <= 0;
        weight_mem[16'h421B] <= 0;
        weight_mem[16'h421C] <= 0;
        weight_mem[16'h421D] <= 0;

        // layer 2 neuron 2
        weight_mem[16'h4400] <= 0;
        weight_mem[16'h4401] <= 0;
        weight_mem[16'h4402] <= 0;
        weight_mem[16'h4403] <= 0;
        weight_mem[16'h4404] <= 0;
        weight_mem[16'h4405] <= 0;
        weight_mem[16'h4406] <= 0;
        weight_mem[16'h4407] <= 0;
        weight_mem[16'h4408] <= 0;
        weight_mem[16'h4409] <= 0;
        weight_mem[16'h440A] <= 0;
        weight_mem[16'h440B] <= 0;
        weight_mem[16'h440C] <= 0;
        weight_mem[16'h440D] <= 0;
        weight_mem[16'h440E] <= 0;
        weight_mem[16'h440F] <= 0;
        weight_mem[16'h4410] <= 0;
        weight_mem[16'h4411] <= 0;
        weight_mem[16'h4412] <= 0;
        weight_mem[16'h4413] <= 0;
        weight_mem[16'h4414] <= 0;
        weight_mem[16'h4415] <= 0;
        weight_mem[16'h4416] <= 0;
        weight_mem[16'h4417] <= 0;
        weight_mem[16'h4418] <= 0;
        weight_mem[16'h4419] <= 0;
        weight_mem[16'h441A] <= 0;
        weight_mem[16'h441B] <= 0;
        weight_mem[16'h441C] <= 0;
        weight_mem[16'h441D] <= 0;

        // layer 2 neuron 3
        weight_mem[16'h4600] <= 0;
        weight_mem[16'h4601] <= 0;
        weight_mem[16'h4602] <= 0;
        weight_mem[16'h4603] <= 0;
        weight_mem[16'h4604] <= 0;
        weight_mem[16'h4605] <= 0;
        weight_mem[16'h4606] <= 0;
        weight_mem[16'h4607] <= 0;
        weight_mem[16'h4608] <= 0;
        weight_mem[16'h4609] <= 0;
        weight_mem[16'h460A] <= 0;
        weight_mem[16'h460B] <= 0;
        weight_mem[16'h460C] <= 0;
        weight_mem[16'h460D] <= 0;
        weight_mem[16'h460E] <= 0;
        weight_mem[16'h460F] <= 0;
        weight_mem[16'h4610] <= 0;
        weight_mem[16'h4611] <= 0;
        weight_mem[16'h4612] <= 0;
        weight_mem[16'h4613] <= 0;
        weight_mem[16'h4614] <= 0;
        weight_mem[16'h4615] <= 0;
        weight_mem[16'h4616] <= 0;
        weight_mem[16'h4617] <= 0;
        weight_mem[16'h4618] <= 0;
        weight_mem[16'h4619] <= 0;
        weight_mem[16'h461A] <= 0;
        weight_mem[16'h461B] <= 0;
        weight_mem[16'h461C] <= 0;
        weight_mem[16'h461D] <= 0;

        // layer 2 neuron 4
        weight_mem[16'h4800] <= 0;
        weight_mem[16'h4801] <= 0;
        weight_mem[16'h4802] <= 0;
        weight_mem[16'h4803] <= 0;
        weight_mem[16'h4804] <= 0;
        weight_mem[16'h4805] <= 0;
        weight_mem[16'h4806] <= 0;
        weight_mem[16'h4807] <= 0;
        weight_mem[16'h4808] <= 0;
        weight_mem[16'h4809] <= 0;
        weight_mem[16'h480A] <= 0;
        weight_mem[16'h480B] <= 0;
        weight_mem[16'h480C] <= 0;
        weight_mem[16'h480D] <= 0;
        weight_mem[16'h480E] <= 0;
        weight_mem[16'h480F] <= 0;
        weight_mem[16'h4810] <= 0;
        weight_mem[16'h4811] <= 0;
        weight_mem[16'h4812] <= 0;
        weight_mem[16'h4813] <= 0;
        weight_mem[16'h4814] <= 0;
        weight_mem[16'h4815] <= 0;
        weight_mem[16'h4816] <= 0;
        weight_mem[16'h4817] <= 0;
        weight_mem[16'h4818] <= 0;
        weight_mem[16'h4819] <= 0;
        weight_mem[16'h481A] <= 0;
        weight_mem[16'h481B] <= 0;
        weight_mem[16'h481C] <= 0;
        weight_mem[16'h481D] <= 0;

        // layer 2 neuron 5
        weight_mem[16'h4A00] <= 0;
        weight_mem[16'h4A01] <= 0;
        weight_mem[16'h4A02] <= 0;
        weight_mem[16'h4A03] <= 0;
        weight_mem[16'h4A04] <= 0;
        weight_mem[16'h4A05] <= 0;
        weight_mem[16'h4A06] <= 0;
        weight_mem[16'h4A07] <= 0;
        weight_mem[16'h4A08] <= 0;
        weight_mem[16'h4A09] <= 0;
        weight_mem[16'h4A0A] <= 0;
        weight_mem[16'h4A0B] <= 0;
        weight_mem[16'h4A0C] <= 0;
        weight_mem[16'h4A0D] <= 0;
        weight_mem[16'h4A0E] <= 0;
        weight_mem[16'h4A0F] <= 0;
        weight_mem[16'h4A10] <= 0;
        weight_mem[16'h4A11] <= 0;
        weight_mem[16'h4A12] <= 0;
        weight_mem[16'h4A13] <= 0;
        weight_mem[16'h4A14] <= 0;
        weight_mem[16'h4A15] <= 0;
        weight_mem[16'h4A16] <= 0;
        weight_mem[16'h4A17] <= 0;
        weight_mem[16'h4A18] <= 0;
        weight_mem[16'h4A19] <= 0;
        weight_mem[16'h4A1A] <= 0;
        weight_mem[16'h4A1B] <= 0;
        weight_mem[16'h4A1C] <= 0;
        weight_mem[16'h4A1D] <= 0;

        // layer 2 neuron 6
        weight_mem[16'h4C00] <= 0;
        weight_mem[16'h4C01] <= 0;
        weight_mem[16'h4C02] <= 0;
        weight_mem[16'h4C03] <= 0;
        weight_mem[16'h4C04] <= 0;
        weight_mem[16'h4C05] <= 0;
        weight_mem[16'h4C06] <= 0;
        weight_mem[16'h4C07] <= 0;
        weight_mem[16'h4C08] <= 0;
        weight_mem[16'h4C09] <= 0;
        weight_mem[16'h4C0A] <= 0;
        weight_mem[16'h4C0B] <= 0;
        weight_mem[16'h4C0C] <= 0;
        weight_mem[16'h4C0D] <= 0;
        weight_mem[16'h4C0E] <= 0;
        weight_mem[16'h4C0F] <= 0;
        weight_mem[16'h4C10] <= 0;
        weight_mem[16'h4C11] <= 0;
        weight_mem[16'h4C12] <= 0;
        weight_mem[16'h4C13] <= 0;
        weight_mem[16'h4C14] <= 0;
        weight_mem[16'h4C15] <= 0;
        weight_mem[16'h4C16] <= 0;
        weight_mem[16'h4C17] <= 0;
        weight_mem[16'h4C18] <= 0;
        weight_mem[16'h4C19] <= 0;
        weight_mem[16'h4C1A] <= 0;
        weight_mem[16'h4C1B] <= 0;
        weight_mem[16'h4C1C] <= 0;
        weight_mem[16'h4C1D] <= 0;

        // layer 2 neuron 7
        weight_mem[16'h4E00] <= 0;
        weight_mem[16'h4E01] <= 0;
        weight_mem[16'h4E02] <= 0;
        weight_mem[16'h4E03] <= 0;
        weight_mem[16'h4E04] <= 0;
        weight_mem[16'h4E05] <= 0;
        weight_mem[16'h4E06] <= 0;
        weight_mem[16'h4E07] <= 0;
        weight_mem[16'h4E08] <= 0;
        weight_mem[16'h4E09] <= 0;
        weight_mem[16'h4E0A] <= 0;
        weight_mem[16'h4E0B] <= 0;
        weight_mem[16'h4E0C] <= 0;
        weight_mem[16'h4E0D] <= 0;
        weight_mem[16'h4E0E] <= 0;
        weight_mem[16'h4E0F] <= 0;
        weight_mem[16'h4E10] <= 0;
        weight_mem[16'h4E11] <= 0;
        weight_mem[16'h4E12] <= 0;
        weight_mem[16'h4E13] <= 0;
        weight_mem[16'h4E14] <= 0;
        weight_mem[16'h4E15] <= 0;
        weight_mem[16'h4E16] <= 0;
        weight_mem[16'h4E17] <= 0;
        weight_mem[16'h4E18] <= 0;
        weight_mem[16'h4E19] <= 0;
        weight_mem[16'h4E1A] <= 0;
        weight_mem[16'h4E1B] <= 0;
        weight_mem[16'h4E1C] <= 0;
        weight_mem[16'h4E1D] <= 0;

        // layer 2 neuron 8
        weight_mem[16'h5000] <= 0;
        weight_mem[16'h5001] <= 0;
        weight_mem[16'h5002] <= 0;
        weight_mem[16'h5003] <= 0;
        weight_mem[16'h5004] <= 0;
        weight_mem[16'h5005] <= 0;
        weight_mem[16'h5006] <= 0;
        weight_mem[16'h5007] <= 0;
        weight_mem[16'h5008] <= 0;
        weight_mem[16'h5009] <= 0;
        weight_mem[16'h500A] <= 0;
        weight_mem[16'h500B] <= 0;
        weight_mem[16'h500C] <= 0;
        weight_mem[16'h500D] <= 0;
        weight_mem[16'h500E] <= 0;
        weight_mem[16'h500F] <= 0;
        weight_mem[16'h5010] <= 0;
        weight_mem[16'h5011] <= 0;
        weight_mem[16'h5012] <= 0;
        weight_mem[16'h5013] <= 0;
        weight_mem[16'h5014] <= 0;
        weight_mem[16'h5015] <= 0;
        weight_mem[16'h5016] <= 0;
        weight_mem[16'h5017] <= 0;
        weight_mem[16'h5018] <= 0;
        weight_mem[16'h5019] <= 0;
        weight_mem[16'h501A] <= 0;
        weight_mem[16'h501B] <= 0;
        weight_mem[16'h501C] <= 0;
        weight_mem[16'h501D] <= 0;

        // layer 2 neuron 9
        weight_mem[16'h5200] <= 0;
        weight_mem[16'h5201] <= 0;
        weight_mem[16'h5202] <= 0;
        weight_mem[16'h5203] <= 0;
        weight_mem[16'h5204] <= 0;
        weight_mem[16'h5205] <= 0;
        weight_mem[16'h5206] <= 0;
        weight_mem[16'h5207] <= 0;
        weight_mem[16'h5208] <= 0;
        weight_mem[16'h5209] <= 0;
        weight_mem[16'h520A] <= 0;
        weight_mem[16'h520B] <= 0;
        weight_mem[16'h520C] <= 0;
        weight_mem[16'h520D] <= 0;
        weight_mem[16'h520E] <= 0;
        weight_mem[16'h520F] <= 0;
        weight_mem[16'h5210] <= 0;
        weight_mem[16'h5211] <= 0;
        weight_mem[16'h5212] <= 0;
        weight_mem[16'h5213] <= 0;
        weight_mem[16'h5214] <= 0;
        weight_mem[16'h5215] <= 0;
        weight_mem[16'h5216] <= 0;
        weight_mem[16'h5217] <= 0;
        weight_mem[16'h5218] <= 0;
        weight_mem[16'h5219] <= 0;
        weight_mem[16'h521A] <= 0;
        weight_mem[16'h521B] <= 0;
        weight_mem[16'h521C] <= 0;
        weight_mem[16'h521D] <= 0;

        // layer 2 neuron 10
        weight_mem[16'h5400] <= 0;
        weight_mem[16'h5401] <= 0;
        weight_mem[16'h5402] <= 0;
        weight_mem[16'h5403] <= 0;
        weight_mem[16'h5404] <= 0;
        weight_mem[16'h5405] <= 0;
        weight_mem[16'h5406] <= 0;
        weight_mem[16'h5407] <= 0;
        weight_mem[16'h5408] <= 0;
        weight_mem[16'h5409] <= 0;
        weight_mem[16'h540A] <= 0;
        weight_mem[16'h540B] <= 0;
        weight_mem[16'h540C] <= 0;
        weight_mem[16'h540D] <= 0;
        weight_mem[16'h540E] <= 0;
        weight_mem[16'h540F] <= 0;
        weight_mem[16'h5410] <= 0;
        weight_mem[16'h5411] <= 0;
        weight_mem[16'h5412] <= 0;
        weight_mem[16'h5413] <= 0;
        weight_mem[16'h5414] <= 0;
        weight_mem[16'h5415] <= 0;
        weight_mem[16'h5416] <= 0;
        weight_mem[16'h5417] <= 0;
        weight_mem[16'h5418] <= 0;
        weight_mem[16'h5419] <= 0;
        weight_mem[16'h541A] <= 0;
        weight_mem[16'h541B] <= 0;
        weight_mem[16'h541C] <= 0;
        weight_mem[16'h541D] <= 0;

        // layer 2 neuron 11
        weight_mem[16'h5600] <= 0;
        weight_mem[16'h5601] <= 0;
        weight_mem[16'h5602] <= 0;
        weight_mem[16'h5603] <= 0;
        weight_mem[16'h5604] <= 0;
        weight_mem[16'h5605] <= 0;
        weight_mem[16'h5606] <= 0;
        weight_mem[16'h5607] <= 0;
        weight_mem[16'h5608] <= 0;
        weight_mem[16'h5609] <= 0;
        weight_mem[16'h560A] <= 0;
        weight_mem[16'h560B] <= 0;
        weight_mem[16'h560C] <= 0;
        weight_mem[16'h560D] <= 0;
        weight_mem[16'h560E] <= 0;
        weight_mem[16'h560F] <= 0;
        weight_mem[16'h5610] <= 0;
        weight_mem[16'h5611] <= 0;
        weight_mem[16'h5612] <= 0;
        weight_mem[16'h5613] <= 0;
        weight_mem[16'h5614] <= 0;
        weight_mem[16'h5615] <= 0;
        weight_mem[16'h5616] <= 0;
        weight_mem[16'h5617] <= 0;
        weight_mem[16'h5618] <= 0;
        weight_mem[16'h5619] <= 0;
        weight_mem[16'h561A] <= 0;
        weight_mem[16'h561B] <= 0;
        weight_mem[16'h561C] <= 0;
        weight_mem[16'h561D] <= 0;

        // layer 2 neuron 12
        weight_mem[16'h5800] <= 0;
        weight_mem[16'h5801] <= 0;
        weight_mem[16'h5802] <= 0;
        weight_mem[16'h5803] <= 0;
        weight_mem[16'h5804] <= 0;
        weight_mem[16'h5805] <= 0;
        weight_mem[16'h5806] <= 0;
        weight_mem[16'h5807] <= 0;
        weight_mem[16'h5808] <= 0;
        weight_mem[16'h5809] <= 0;
        weight_mem[16'h580A] <= 0;
        weight_mem[16'h580B] <= 0;
        weight_mem[16'h580C] <= 0;
        weight_mem[16'h580D] <= 0;
        weight_mem[16'h580E] <= 0;
        weight_mem[16'h580F] <= 0;
        weight_mem[16'h5810] <= 0;
        weight_mem[16'h5811] <= 0;
        weight_mem[16'h5812] <= 0;
        weight_mem[16'h5813] <= 0;
        weight_mem[16'h5814] <= 0;
        weight_mem[16'h5815] <= 0;
        weight_mem[16'h5816] <= 0;
        weight_mem[16'h5817] <= 0;
        weight_mem[16'h5818] <= 0;
        weight_mem[16'h5819] <= 0;
        weight_mem[16'h581A] <= 0;
        weight_mem[16'h581B] <= 0;
        weight_mem[16'h581C] <= 0;
        weight_mem[16'h581D] <= 0;

        // layer 2 neuron 13
        weight_mem[16'h5A00] <= 0;
        weight_mem[16'h5A01] <= 0;
        weight_mem[16'h5A02] <= 0;
        weight_mem[16'h5A03] <= 0;
        weight_mem[16'h5A04] <= 0;
        weight_mem[16'h5A05] <= 0;
        weight_mem[16'h5A06] <= 0;
        weight_mem[16'h5A07] <= 0;
        weight_mem[16'h5A08] <= 0;
        weight_mem[16'h5A09] <= 0;
        weight_mem[16'h5A0A] <= 0;
        weight_mem[16'h5A0B] <= 0;
        weight_mem[16'h5A0C] <= 0;
        weight_mem[16'h5A0D] <= 0;
        weight_mem[16'h5A0E] <= 0;
        weight_mem[16'h5A0F] <= 0;
        weight_mem[16'h5A10] <= 0;
        weight_mem[16'h5A11] <= 0;
        weight_mem[16'h5A12] <= 0;
        weight_mem[16'h5A13] <= 0;
        weight_mem[16'h5A14] <= 0;
        weight_mem[16'h5A15] <= 0;
        weight_mem[16'h5A16] <= 0;
        weight_mem[16'h5A17] <= 0;
        weight_mem[16'h5A18] <= 0;
        weight_mem[16'h5A19] <= 0;
        weight_mem[16'h5A1A] <= 0;
        weight_mem[16'h5A1B] <= 0;
        weight_mem[16'h5A1C] <= 0;
        weight_mem[16'h5A1D] <= 0;

        // layer 2 neuron 14
        weight_mem[16'h5C00] <= 0;
        weight_mem[16'h5C01] <= 0;
        weight_mem[16'h5C02] <= 0;
        weight_mem[16'h5C03] <= 0;
        weight_mem[16'h5C04] <= 0;
        weight_mem[16'h5C05] <= 0;
        weight_mem[16'h5C06] <= 0;
        weight_mem[16'h5C07] <= 0;
        weight_mem[16'h5C08] <= 0;
        weight_mem[16'h5C09] <= 0;
        weight_mem[16'h5C0A] <= 0;
        weight_mem[16'h5C0B] <= 0;
        weight_mem[16'h5C0C] <= 0;
        weight_mem[16'h5C0D] <= 0;
        weight_mem[16'h5C0E] <= 0;
        weight_mem[16'h5C0F] <= 0;
        weight_mem[16'h5C10] <= 0;
        weight_mem[16'h5C11] <= 0;
        weight_mem[16'h5C12] <= 0;
        weight_mem[16'h5C13] <= 0;
        weight_mem[16'h5C14] <= 0;
        weight_mem[16'h5C15] <= 0;
        weight_mem[16'h5C16] <= 0;
        weight_mem[16'h5C17] <= 0;
        weight_mem[16'h5C18] <= 0;
        weight_mem[16'h5C19] <= 0;
        weight_mem[16'h5C1A] <= 0;
        weight_mem[16'h5C1B] <= 0;
        weight_mem[16'h5C1C] <= 0;
        weight_mem[16'h5C1D] <= 0;

        // layer 2 neuron 15
        weight_mem[16'h5E00] <= 0;
        weight_mem[16'h5E01] <= 0;
        weight_mem[16'h5E02] <= 0;
        weight_mem[16'h5E03] <= 0;
        weight_mem[16'h5E04] <= 0;
        weight_mem[16'h5E05] <= 0;
        weight_mem[16'h5E06] <= 0;
        weight_mem[16'h5E07] <= 0;
        weight_mem[16'h5E08] <= 0;
        weight_mem[16'h5E09] <= 0;
        weight_mem[16'h5E0A] <= 0;
        weight_mem[16'h5E0B] <= 0;
        weight_mem[16'h5E0C] <= 0;
        weight_mem[16'h5E0D] <= 0;
        weight_mem[16'h5E0E] <= 0;
        weight_mem[16'h5E0F] <= 0;
        weight_mem[16'h5E10] <= 0;
        weight_mem[16'h5E11] <= 0;
        weight_mem[16'h5E12] <= 0;
        weight_mem[16'h5E13] <= 0;
        weight_mem[16'h5E14] <= 0;
        weight_mem[16'h5E15] <= 0;
        weight_mem[16'h5E16] <= 0;
        weight_mem[16'h5E17] <= 0;
        weight_mem[16'h5E18] <= 0;
        weight_mem[16'h5E19] <= 0;
        weight_mem[16'h5E1A] <= 0;
        weight_mem[16'h5E1B] <= 0;
        weight_mem[16'h5E1C] <= 0;
        weight_mem[16'h5E1D] <= 0;

        // layer 3 neuron 0
        weight_mem[16'h8000] <= 0;
        weight_mem[16'h8001] <= 0;
        weight_mem[16'h8002] <= 0;
        weight_mem[16'h8003] <= 0;
        weight_mem[16'h8004] <= 0;
        weight_mem[16'h8005] <= 0;
        weight_mem[16'h8006] <= 0;
        weight_mem[16'h8007] <= 0;
        weight_mem[16'h8008] <= 0;
        weight_mem[16'h8009] <= 0;
        weight_mem[16'h800A] <= 0;
        weight_mem[16'h800B] <= 0;
        weight_mem[16'h800C] <= 0;
        weight_mem[16'h800D] <= 0;
        weight_mem[16'h800E] <= 0;
        weight_mem[16'h800F] <= 0;

        // layer 3 neuron 1
        weight_mem[16'h8200] <= 1;
        weight_mem[16'h8201] <= 0;
        weight_mem[16'h8202] <= 0;
        weight_mem[16'h8203] <= 0;
        weight_mem[16'h8204] <= 0;
        weight_mem[16'h8205] <= 0;
        weight_mem[16'h8206] <= 0;
        weight_mem[16'h8207] <= 0;
        weight_mem[16'h8208] <= 0;
        weight_mem[16'h8209] <= 0;
        weight_mem[16'h820A] <= 0;
        weight_mem[16'h820B] <= 0;
        weight_mem[16'h820C] <= 0;
        weight_mem[16'h820D] <= 0;
        weight_mem[16'h820E] <= 0;
        weight_mem[16'h820F] <= 0;

        // layer 3 neuron 2
        weight_mem[16'h8400] <= 2;
        weight_mem[16'h8401] <= 0;
        weight_mem[16'h8402] <= 0;
        weight_mem[16'h8403] <= 0;
        weight_mem[16'h8404] <= 0;
        weight_mem[16'h8405] <= 0;
        weight_mem[16'h8406] <= 0;
        weight_mem[16'h8407] <= 0;
        weight_mem[16'h8408] <= 0;
        weight_mem[16'h8409] <= 0;
        weight_mem[16'h840A] <= 0;
        weight_mem[16'h840B] <= 0;
        weight_mem[16'h840C] <= 0;
        weight_mem[16'h840D] <= 0;
        weight_mem[16'h840E] <= 0;
        weight_mem[16'h840F] <= 0;

        // layer 3 neuron 3
        weight_mem[16'h8600] <= 3;
        weight_mem[16'h8601] <= 0;
        weight_mem[16'h8602] <= 0;
        weight_mem[16'h8603] <= 0;
        weight_mem[16'h8604] <= 0;
        weight_mem[16'h8605] <= 0;
        weight_mem[16'h8606] <= 0;
        weight_mem[16'h8607] <= 0;
        weight_mem[16'h8608] <= 0;
        weight_mem[16'h8609] <= 0;
        weight_mem[16'h860A] <= 0;
        weight_mem[16'h860B] <= 0;
        weight_mem[16'h860C] <= 0;
        weight_mem[16'h860D] <= 0;
        weight_mem[16'h860E] <= 0;
        weight_mem[16'h860F] <= 0;

        // layer 3 neuron 4
        weight_mem[16'h8800] <= 4;
        weight_mem[16'h8801] <= 0;
        weight_mem[16'h8802] <= 0;
        weight_mem[16'h8803] <= 0;
        weight_mem[16'h8804] <= 0;
        weight_mem[16'h8805] <= 0;
        weight_mem[16'h8806] <= 0;
        weight_mem[16'h8807] <= 0;
        weight_mem[16'h8808] <= 0;
        weight_mem[16'h8809] <= 0;
        weight_mem[16'h880A] <= 0;
        weight_mem[16'h880B] <= 0;
        weight_mem[16'h880C] <= 0;
        weight_mem[16'h880D] <= 0;
        weight_mem[16'h880E] <= 0;
        weight_mem[16'h880F] <= 0;

        // layer 3 neuron 5
        weight_mem[16'h8A00] <= 5;
        weight_mem[16'h8A01] <= 0;
        weight_mem[16'h8A02] <= 0;
        weight_mem[16'h8A03] <= 0;
        weight_mem[16'h8A04] <= 0;
        weight_mem[16'h8A05] <= 0;
        weight_mem[16'h8A06] <= 0;
        weight_mem[16'h8A07] <= 0;
        weight_mem[16'h8A08] <= 0;
        weight_mem[16'h8A09] <= 0;
        weight_mem[16'h8A0A] <= 0;
        weight_mem[16'h8A0B] <= 0;
        weight_mem[16'h8A0C] <= 0;
        weight_mem[16'h8A0D] <= 0;
        weight_mem[16'h8A0E] <= 0;
        weight_mem[16'h8A0F] <= 0;

        // layer 3 neuron 6
        weight_mem[16'h8C00] <= 6;
        weight_mem[16'h8C01] <= 0;
        weight_mem[16'h8C02] <= 0;
        weight_mem[16'h8C03] <= 0;
        weight_mem[16'h8C04] <= 0;
        weight_mem[16'h8C05] <= 0;
        weight_mem[16'h8C06] <= 0;
        weight_mem[16'h8C07] <= 0;
        weight_mem[16'h8C08] <= 0;
        weight_mem[16'h8C09] <= 0;
        weight_mem[16'h8C0A] <= 0;
        weight_mem[16'h8C0B] <= 0;
        weight_mem[16'h8C0C] <= 0;
        weight_mem[16'h8C0D] <= 0;
        weight_mem[16'h8C0E] <= 0;
        weight_mem[16'h8C0F] <= 0;

        // layer 3 neuron 7
        weight_mem[16'h8E00] <= 7;
        weight_mem[16'h8E01] <= 0;
        weight_mem[16'h8E02] <= 0;
        weight_mem[16'h8E03] <= 0;
        weight_mem[16'h8E04] <= 0;
        weight_mem[16'h8E05] <= 0;
        weight_mem[16'h8E06] <= 0;
        weight_mem[16'h8E07] <= 0;
        weight_mem[16'h8E08] <= 0;
        weight_mem[16'h8E09] <= 0;
        weight_mem[16'h8E0A] <= 0;
        weight_mem[16'h8E0B] <= 0;
        weight_mem[16'h8E0C] <= 0;
        weight_mem[16'h8E0D] <= 0;
        weight_mem[16'h8E0E] <= 0;
        weight_mem[16'h8E0F] <= 0;

        // layer 3 neuron 8
        weight_mem[16'h9000] <= 8;
        weight_mem[16'h9001] <= 0;
        weight_mem[16'h9002] <= 0;
        weight_mem[16'h9003] <= 0;
        weight_mem[16'h9004] <= 0;
        weight_mem[16'h9005] <= 0;
        weight_mem[16'h9006] <= 0;
        weight_mem[16'h9007] <= 0;
        weight_mem[16'h9008] <= 0;
        weight_mem[16'h9009] <= 0;
        weight_mem[16'h900A] <= 0;
        weight_mem[16'h900B] <= 0;
        weight_mem[16'h900C] <= 0;
        weight_mem[16'h900D] <= 0;
        weight_mem[16'h900E] <= 0;
        weight_mem[16'h900F] <= 0;

        // layer 3 neuron 9
        weight_mem[16'h9200] <= 9;
        weight_mem[16'h9201] <= 0;
        weight_mem[16'h9202] <= 0;
        weight_mem[16'h9203] <= 0;
        weight_mem[16'h9204] <= 0;
        weight_mem[16'h9205] <= 0;
        weight_mem[16'h9206] <= 0;
        weight_mem[16'h9207] <= 0;
        weight_mem[16'h9208] <= 0;
        weight_mem[16'h9209] <= 0;
        weight_mem[16'h920A] <= 0;
        weight_mem[16'h920B] <= 0;
        weight_mem[16'h920C] <= 0;
        weight_mem[16'h920D] <= 0;
        weight_mem[16'h920E] <= 0;
        weight_mem[16'h920F] <= 0;

    end

    always @(posedge clk) begin
        if (reset) begin
            weight_val <= 0;
        end else begin 
            weight_val <= weight_mem[input_addr];
        end
    end

endmodule

