module neuron_mem
    (
        input wire clk, 
        input wire reset,
        input wire write_enable,
        input wire [11:0] input_addr,
        input wire signed [15:0] data,
        input wire [11:0] output_addr,
        output reg signed [15:0] neuron_val
    );

    // 2^12 (size of neuron address) requires 4096 addresses
    reg signed [15:0] neuron_mem[0:4095];

    // initializing input layer
    initial begin
        neuron_mem[0] <= 1;
        neuron_mem[1] <= 0;
        neuron_mem[2] <= 0;
        neuron_mem[3] <= 0;
        neuron_mem[4] <= 0;
        neuron_mem[5] <= 0;
        neuron_mem[6] <= 0;
        neuron_mem[7] <= 0;
        neuron_mem[8] <= 0;
        neuron_mem[9] <= 0;
        neuron_mem[10] <= 0;
        neuron_mem[11] <= 0;
        neuron_mem[12] <= 0;
        neuron_mem[13] <= 0;
        neuron_mem[14] <= 0;
        neuron_mem[15] <= 0;
        neuron_mem[16] <= 0;
        neuron_mem[17] <= 0;
        neuron_mem[18] <= 0;
        neuron_mem[19] <= 0;
        neuron_mem[20] <= 0;
        neuron_mem[21] <= 0;
        neuron_mem[22] <= 0;
        neuron_mem[23] <= 0;
        neuron_mem[24] <= 0;
        neuron_mem[25] <= 0;
        neuron_mem[26] <= 0;
        neuron_mem[27] <= 0;
        neuron_mem[28] <= 0;
        neuron_mem[29] <= 0;
        neuron_mem[30] <= 0;
        neuron_mem[31] <= 0;
        neuron_mem[32] <= 0;
        neuron_mem[33] <= 0;
        neuron_mem[34] <= 0;
        neuron_mem[35] <= 0;
        neuron_mem[36] <= 0;
        neuron_mem[37] <= 0;
        neuron_mem[38] <= 0;
        neuron_mem[39] <= 0;
        neuron_mem[40] <= 0;
        neuron_mem[41] <= 0;
        neuron_mem[42] <= 0;
        neuron_mem[43] <= 0;
        neuron_mem[44] <= 0;
        neuron_mem[45] <= 0;
        neuron_mem[46] <= 0;
        neuron_mem[47] <= 0;
        neuron_mem[48] <= 0;
        neuron_mem[49] <= 0;
        neuron_mem[50] <= 0;
        neuron_mem[51] <= 0;
        neuron_mem[52] <= 0;
        neuron_mem[53] <= 0;
        neuron_mem[54] <= 0;
        neuron_mem[55] <= 0;
        neuron_mem[56] <= 0;
        neuron_mem[57] <= 0;
        neuron_mem[58] <= 0;
        neuron_mem[59] <= 0;
        neuron_mem[60] <= 0;
        neuron_mem[61] <= 0;
        neuron_mem[62] <= 0;
        neuron_mem[63] <= 0;
        neuron_mem[64] <= 0;
        neuron_mem[65] <= 0;
        neuron_mem[66] <= 0;
        neuron_mem[67] <= 0;
        neuron_mem[68] <= 0;
        neuron_mem[69] <= 0;
        neuron_mem[70] <= 0;
        neuron_mem[71] <= 0;
        neuron_mem[72] <= 0;
        neuron_mem[73] <= 0;
        neuron_mem[74] <= 0;
        neuron_mem[75] <= 0;
        neuron_mem[76] <= 0;
        neuron_mem[77] <= 0;
        neuron_mem[78] <= 0;
        neuron_mem[79] <= 0;
        neuron_mem[80] <= 0;
        neuron_mem[81] <= 0;
        neuron_mem[82] <= 0;
        neuron_mem[83] <= 0;
        neuron_mem[84] <= 0;
        neuron_mem[85] <= 0;
        neuron_mem[86] <= 0;
        neuron_mem[87] <= 0;
        neuron_mem[88] <= 0;
        neuron_mem[89] <= 0;
        neuron_mem[90] <= 0;
        neuron_mem[91] <= 0;
        neuron_mem[92] <= 0;
        neuron_mem[93] <= 0;
        neuron_mem[94] <= 0;
        neuron_mem[95] <= 0;
        neuron_mem[96] <= 0;
        neuron_mem[97] <= 0;
        neuron_mem[98] <= 0;
        neuron_mem[99] <= 0;
        neuron_mem[100] <= 0;
        neuron_mem[101] <= 0;
        neuron_mem[102] <= 0;
        neuron_mem[103] <= 0;
        neuron_mem[104] <= 0;
        neuron_mem[105] <= 0;
        neuron_mem[106] <= 0;
        neuron_mem[107] <= 0;
        neuron_mem[108] <= 0;
        neuron_mem[109] <= 0;
        neuron_mem[110] <= 0;
        neuron_mem[111] <= 0;
        neuron_mem[112] <= 0;
        neuron_mem[113] <= 0;
        neuron_mem[114] <= 0;
        neuron_mem[115] <= 0;
        neuron_mem[116] <= 0;
        neuron_mem[117] <= 0;
        neuron_mem[118] <= 0;
        neuron_mem[119] <= 0;
        neuron_mem[120] <= 0;
        neuron_mem[121] <= 0;
        neuron_mem[122] <= 0;
        neuron_mem[123] <= 0;
        neuron_mem[124] <= 0;
        neuron_mem[125] <= 0;
        neuron_mem[126] <= 0;
        neuron_mem[127] <= 0;
        neuron_mem[128] <= 0;
        neuron_mem[129] <= 0;
        neuron_mem[130] <= 0;
        neuron_mem[131] <= 0;
        neuron_mem[132] <= 0;
        neuron_mem[133] <= 0;
        neuron_mem[134] <= 0;
        neuron_mem[135] <= 0;
        neuron_mem[136] <= 0;
        neuron_mem[137] <= 0;
        neuron_mem[138] <= 0;
        neuron_mem[139] <= 0;
        neuron_mem[140] <= 0;
        neuron_mem[141] <= 0;
        neuron_mem[142] <= 0;
        neuron_mem[143] <= 0;
        neuron_mem[144] <= 0;
        neuron_mem[145] <= 0;
        neuron_mem[146] <= 0;
        neuron_mem[147] <= 0;
        neuron_mem[148] <= 0;
        neuron_mem[149] <= 0;
        neuron_mem[150] <= 0;
        neuron_mem[151] <= 0;
        neuron_mem[152] <= 0;
        neuron_mem[153] <= 0;
        neuron_mem[154] <= 0;
        neuron_mem[155] <= 0;
        neuron_mem[156] <= 0;
        neuron_mem[157] <= 0;
        neuron_mem[158] <= 0;
        neuron_mem[159] <= 0;
        neuron_mem[160] <= 0;
        neuron_mem[161] <= 0;
        neuron_mem[162] <= 0;
        neuron_mem[163] <= 0;
        neuron_mem[164] <= 0;
        neuron_mem[165] <= 0;
        neuron_mem[166] <= 0;
        neuron_mem[167] <= 0;
        neuron_mem[168] <= 0;
        neuron_mem[169] <= 0;
        neuron_mem[170] <= 0;
        neuron_mem[171] <= 0;
        neuron_mem[172] <= 0;
        neuron_mem[173] <= 0;
        neuron_mem[174] <= 0;
        neuron_mem[175] <= 0;
        neuron_mem[176] <= 0;
        neuron_mem[177] <= 0;
        neuron_mem[178] <= 0;
        neuron_mem[179] <= 0;
        neuron_mem[180] <= 0;
        neuron_mem[181] <= 0;
        neuron_mem[182] <= 0;
        neuron_mem[183] <= 0;
        neuron_mem[184] <= 0;
        neuron_mem[185] <= 0;
        neuron_mem[186] <= 0;
        neuron_mem[187] <= 0;
        neuron_mem[188] <= 0;
        neuron_mem[189] <= 0;
        neuron_mem[190] <= 0;
        neuron_mem[191] <= 0;
        neuron_mem[192] <= 0;
        neuron_mem[193] <= 0;
        neuron_mem[194] <= 0;
        neuron_mem[195] <= 0;
        neuron_mem[196] <= 0;
        neuron_mem[197] <= 0;
        neuron_mem[198] <= 0;
        neuron_mem[199] <= 0;
        neuron_mem[200] <= 0;
        neuron_mem[201] <= 0;
        neuron_mem[202] <= 0;
        neuron_mem[203] <= 0;
        neuron_mem[204] <= 0;
        neuron_mem[205] <= 0;
        neuron_mem[206] <= 0;
        neuron_mem[207] <= 0;
        neuron_mem[208] <= 0;
        neuron_mem[209] <= 0;
        neuron_mem[210] <= 0;
        neuron_mem[211] <= 0;
        neuron_mem[212] <= 0;
        neuron_mem[213] <= 0;
        neuron_mem[214] <= 0;
        neuron_mem[215] <= 0;
        neuron_mem[216] <= 0;
        neuron_mem[217] <= 0;
        neuron_mem[218] <= 0;
        neuron_mem[219] <= 0;
        neuron_mem[220] <= 0;
        neuron_mem[221] <= 0;
        neuron_mem[222] <= 0;
        neuron_mem[223] <= 0;
        neuron_mem[224] <= 0;
        neuron_mem[225] <= 0;
        neuron_mem[226] <= 0;
        neuron_mem[227] <= 0;
        neuron_mem[228] <= 0;
        neuron_mem[229] <= 0;
        neuron_mem[230] <= 0;
        neuron_mem[231] <= 0;
        neuron_mem[232] <= 0;
        neuron_mem[233] <= 0;
        neuron_mem[234] <= 0;
        neuron_mem[235] <= 0;
        neuron_mem[236] <= 0;
        neuron_mem[237] <= 0;
        neuron_mem[238] <= 0;
        neuron_mem[239] <= 0;
        neuron_mem[240] <= 0;
        neuron_mem[241] <= 0;
        neuron_mem[242] <= 0;
        neuron_mem[243] <= 0;
        neuron_mem[244] <= 0;
        neuron_mem[245] <= 0;
        neuron_mem[246] <= 0;
        neuron_mem[247] <= 0;
        neuron_mem[248] <= 0;
        neuron_mem[249] <= 0;
        neuron_mem[250] <= 0;
        neuron_mem[251] <= 0;
        neuron_mem[252] <= 0;
        neuron_mem[253] <= 0;
        neuron_mem[254] <= 0;
        neuron_mem[255] <= 0;
        neuron_mem[256] <= 0;
        neuron_mem[257] <= 0;
        neuron_mem[258] <= 0;
        neuron_mem[259] <= 0;
        neuron_mem[260] <= 0;
        neuron_mem[261] <= 0;
        neuron_mem[262] <= 0;
        neuron_mem[263] <= 0;
        neuron_mem[264] <= 0;
        neuron_mem[265] <= 0;
        neuron_mem[266] <= 0;
        neuron_mem[267] <= 0;
        neuron_mem[268] <= 0;
        neuron_mem[269] <= 0;
        neuron_mem[270] <= 0;
        neuron_mem[271] <= 0;
        neuron_mem[272] <= 0;
        neuron_mem[273] <= 0;
        neuron_mem[274] <= 0;
        neuron_mem[275] <= 0;
        neuron_mem[276] <= 0;
        neuron_mem[277] <= 0;
        neuron_mem[278] <= 0;
        neuron_mem[279] <= 0;
        neuron_mem[280] <= 0;
        neuron_mem[281] <= 0;
        neuron_mem[282] <= 0;
        neuron_mem[283] <= 0;
        neuron_mem[284] <= 0;
        neuron_mem[285] <= 0;
        neuron_mem[286] <= 0;
        neuron_mem[287] <= 0;
        neuron_mem[288] <= 0;
        neuron_mem[289] <= 0;
        neuron_mem[290] <= 0;
        neuron_mem[291] <= 0;
        neuron_mem[292] <= 0;
        neuron_mem[293] <= 0;
        neuron_mem[294] <= 0;
        neuron_mem[295] <= 0;
        neuron_mem[296] <= 0;
        neuron_mem[297] <= 0;
        neuron_mem[298] <= 0;
        neuron_mem[299] <= 0;
        neuron_mem[300] <= 0;
        neuron_mem[301] <= 0;
        neuron_mem[302] <= 0;
        neuron_mem[303] <= 0;
        neuron_mem[304] <= 0;
        neuron_mem[305] <= 0;
        neuron_mem[306] <= 0;
        neuron_mem[307] <= 0;
        neuron_mem[308] <= 0;
        neuron_mem[309] <= 0;
        neuron_mem[310] <= 0;
        neuron_mem[311] <= 0;
        neuron_mem[312] <= 0;
        neuron_mem[313] <= 0;
        neuron_mem[314] <= 0;
        neuron_mem[315] <= 0;
        neuron_mem[316] <= 0;
        neuron_mem[317] <= 0;
        neuron_mem[318] <= 0;
        neuron_mem[319] <= 0;
        neuron_mem[320] <= 0;
        neuron_mem[321] <= 0;
        neuron_mem[322] <= 0;
        neuron_mem[323] <= 0;
        neuron_mem[324] <= 0;
        neuron_mem[325] <= 0;
        neuron_mem[326] <= 0;
        neuron_mem[327] <= 0;
        neuron_mem[328] <= 0;
        neuron_mem[329] <= 0;
        neuron_mem[330] <= 0;
        neuron_mem[331] <= 0;
        neuron_mem[332] <= 0;
        neuron_mem[333] <= 0;
        neuron_mem[334] <= 0;
        neuron_mem[335] <= 0;
        neuron_mem[336] <= 0;
        neuron_mem[337] <= 0;
        neuron_mem[338] <= 0;
        neuron_mem[339] <= 0;
        neuron_mem[340] <= 0;
        neuron_mem[341] <= 0;
        neuron_mem[342] <= 0;
        neuron_mem[343] <= 0;
        neuron_mem[344] <= 0;
        neuron_mem[345] <= 0;
        neuron_mem[346] <= 0;
        neuron_mem[347] <= 0;
        neuron_mem[348] <= 0;
        neuron_mem[349] <= 0;
        neuron_mem[350] <= 0;
        neuron_mem[351] <= 0;
        neuron_mem[352] <= 0;
        neuron_mem[353] <= 0;
        neuron_mem[354] <= 0;
        neuron_mem[355] <= 0;
        neuron_mem[356] <= 0;
        neuron_mem[357] <= 0;
        neuron_mem[358] <= 0;
        neuron_mem[359] <= 0;
        neuron_mem[360] <= 0;
        neuron_mem[361] <= 0;
        neuron_mem[362] <= 0;
        neuron_mem[363] <= 0;
        neuron_mem[364] <= 0;
        neuron_mem[365] <= 0;
        neuron_mem[366] <= 0;
        neuron_mem[367] <= 0;
        neuron_mem[368] <= 0;
        neuron_mem[369] <= 0;
        neuron_mem[370] <= 0;
        neuron_mem[371] <= 0;
        neuron_mem[372] <= 0;
        neuron_mem[373] <= 0;
        neuron_mem[374] <= 0;
        neuron_mem[375] <= 0;
        neuron_mem[376] <= 0;
        neuron_mem[377] <= 0;
        neuron_mem[378] <= 0;
        neuron_mem[379] <= 0;
        neuron_mem[380] <= 0;
        neuron_mem[381] <= 0;
        neuron_mem[382] <= 0;
        neuron_mem[383] <= 0;
        neuron_mem[384] <= 0;
        neuron_mem[385] <= 0;
        neuron_mem[386] <= 0;
        neuron_mem[387] <= 0;
        neuron_mem[388] <= 0;
        neuron_mem[389] <= 0;
        neuron_mem[390] <= 0;
        neuron_mem[391] <= 0;
        neuron_mem[392] <= 0;
        neuron_mem[393] <= 0;
        neuron_mem[394] <= 0;
        neuron_mem[395] <= 0;
        neuron_mem[396] <= 0;
        neuron_mem[397] <= 0;
        neuron_mem[398] <= 0;
        neuron_mem[399] <= 0;
        neuron_mem[400] <= 0;
        neuron_mem[401] <= 0;
        neuron_mem[402] <= 0;
        neuron_mem[403] <= 0;
        neuron_mem[404] <= 0;
        neuron_mem[405] <= 0;
        neuron_mem[406] <= 0;
        neuron_mem[407] <= 0;
        neuron_mem[408] <= 0;
        neuron_mem[409] <= 0;
        neuron_mem[410] <= 0;
        neuron_mem[411] <= 0;
        neuron_mem[412] <= 0;
        neuron_mem[413] <= 0;
        neuron_mem[414] <= 0;
        neuron_mem[415] <= 0;
        neuron_mem[416] <= 0;
        neuron_mem[417] <= 0;
        neuron_mem[418] <= 0;
        neuron_mem[419] <= 0;
        neuron_mem[420] <= 0;
        neuron_mem[421] <= 0;
        neuron_mem[422] <= 0;
        neuron_mem[423] <= 0;
        neuron_mem[424] <= 0;
        neuron_mem[425] <= 0;
        neuron_mem[426] <= 0;
        neuron_mem[427] <= 0;
        neuron_mem[428] <= 0;
        neuron_mem[429] <= 0;
        neuron_mem[430] <= 0;
        neuron_mem[431] <= 0;
    end

    always @(posedge clk) begin
        if (reset) begin
            neuron_val <= 0;
        end else begin 
            if (input_addr == output_addr && write_enable) begin
                neuron_val <= data;
            end else begin
                neuron_val <= neuron_mem[input_addr];
            end 

            if (write_enable) begin
                neuron_mem[output_addr] <= data;
            end
        end
    end

endmodule
