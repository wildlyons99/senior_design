module weight_mem
    (
        input wire clk, 
        input wire reset,
        input wire [15:0] input_addr,
        output reg signed [7:0] weight_val
    );

    // 2^16 (size of neuron address) requires 65536 addresses
    reg signed [7:0] weight_mem[0:65535];

    // initializing input layer
    initial begin
        // layer 1 neuron 0
        weight_mem[16'h0000] <= 254;
        weight_mem[16'h0001] <= 3;
        weight_mem[16'h0002] <= 247;
        weight_mem[16'h0003] <= 247;
        weight_mem[16'h0004] <= 243;
        weight_mem[16'h0005] <= 7;
        weight_mem[16'h0006] <= 253;
        weight_mem[16'h0007] <= 245;
        weight_mem[16'h0008] <= 248;
        weight_mem[16'h0009] <= 0;
        weight_mem[16'h000A] <= 241;
        weight_mem[16'h000B] <= 241;
        weight_mem[16'h000C] <= 249;
        weight_mem[16'h000D] <= 251;
        weight_mem[16'h000E] <= 249;
        weight_mem[16'h000F] <= 245;
        weight_mem[16'h0010] <= 252;
        weight_mem[16'h0011] <= 250;
        weight_mem[16'h0012] <= 248;
        weight_mem[16'h0013] <= 2;
        weight_mem[16'h0014] <= 4;
        weight_mem[16'h0015] <= 248;
        weight_mem[16'h0016] <= 0;
        weight_mem[16'h0017] <= 252;
        weight_mem[16'h0018] <= 247;
        weight_mem[16'h0019] <= 247;
        weight_mem[16'h001A] <= 4;
        weight_mem[16'h001B] <= 254;
        weight_mem[16'h001C] <= 254;
        weight_mem[16'h001D] <= 253;
        weight_mem[16'h001E] <= 3;
        weight_mem[16'h001F] <= 0;
        weight_mem[16'h0020] <= 246;
        weight_mem[16'h0021] <= 241;
        weight_mem[16'h0022] <= 241;
        weight_mem[16'h0023] <= 242;
        weight_mem[16'h0024] <= 3;
        weight_mem[16'h0025] <= 248;
        weight_mem[16'h0026] <= 248;
        weight_mem[16'h0027] <= 7;
        weight_mem[16'h0028] <= 253;
        weight_mem[16'h0029] <= 244;
        weight_mem[16'h002A] <= 242;
        weight_mem[16'h002B] <= 246;
        weight_mem[16'h002C] <= 0;
        weight_mem[16'h002D] <= 241;
        weight_mem[16'h002E] <= 5;
        weight_mem[16'h002F] <= 245;
        weight_mem[16'h0030] <= 249;
        weight_mem[16'h0031] <= 244;
        weight_mem[16'h0032] <= 253;
        weight_mem[16'h0033] <= 5;
        weight_mem[16'h0034] <= 1;
        weight_mem[16'h0035] <= 4;
        weight_mem[16'h0036] <= 252;
        weight_mem[16'h0037] <= 1;
        weight_mem[16'h0038] <= 251;
        weight_mem[16'h0039] <= 0;
        weight_mem[16'h003A] <= 0;
        weight_mem[16'h003B] <= 245;
        weight_mem[16'h003C] <= 1;
        weight_mem[16'h003D] <= 20;
        weight_mem[16'h003E] <= 17;
        weight_mem[16'h003F] <= 24;
        weight_mem[16'h0040] <= 11;
        weight_mem[16'h0041] <= 13;
        weight_mem[16'h0042] <= 10;
        weight_mem[16'h0043] <= 7;
        weight_mem[16'h0044] <= 241;
        weight_mem[16'h0045] <= 241;
        weight_mem[16'h0046] <= 251;
        weight_mem[16'h0047] <= 246;
        weight_mem[16'h0048] <= 5;
        weight_mem[16'h0049] <= 255;
        weight_mem[16'h004A] <= 3;
        weight_mem[16'h004B] <= 252;
        weight_mem[16'h004C] <= 251;
        weight_mem[16'h004D] <= 253;
        weight_mem[16'h004E] <= 230;
        weight_mem[16'h004F] <= 233;
        weight_mem[16'h0050] <= 229;
        weight_mem[16'h0051] <= 2;
        weight_mem[16'h0052] <= 5;
        weight_mem[16'h0053] <= 16;
        weight_mem[16'h0054] <= 46;
        weight_mem[16'h0055] <= 45;
        weight_mem[16'h0056] <= 64;
        weight_mem[16'h0057] <= 44;
        weight_mem[16'h0058] <= 51;
        weight_mem[16'h0059] <= 29;
        weight_mem[16'h005A] <= 22;
        weight_mem[16'h005B] <= 15;
        weight_mem[16'h005C] <= 249;
        weight_mem[16'h005D] <= 254;
        weight_mem[16'h005E] <= 2;
        weight_mem[16'h005F] <= 245;
        weight_mem[16'h0060] <= 0;
        weight_mem[16'h0061] <= 253;
        weight_mem[16'h0062] <= 247;
        weight_mem[16'h0063] <= 238;
        weight_mem[16'h0064] <= 246;
        weight_mem[16'h0065] <= 235;
        weight_mem[16'h0066] <= 233;
        weight_mem[16'h0067] <= 232;
        weight_mem[16'h0068] <= 250;
        weight_mem[16'h0069] <= 250;
        weight_mem[16'h006A] <= 9;
        weight_mem[16'h006B] <= 10;
        weight_mem[16'h006C] <= 27;
        weight_mem[16'h006D] <= 45;
        weight_mem[16'h006E] <= 27;
        weight_mem[16'h006F] <= 51;
        weight_mem[16'h0070] <= 35;
        weight_mem[16'h0071] <= 40;
        weight_mem[16'h0072] <= 16;
        weight_mem[16'h0073] <= 15;
        weight_mem[16'h0074] <= 18;
        weight_mem[16'h0075] <= 18;
        weight_mem[16'h0076] <= 13;
        weight_mem[16'h0077] <= 244;
        weight_mem[16'h0078] <= 3;
        weight_mem[16'h0079] <= 251;
        weight_mem[16'h007A] <= 253;
        weight_mem[16'h007B] <= 230;
        weight_mem[16'h007C] <= 228;
        weight_mem[16'h007D] <= 235;
        weight_mem[16'h007E] <= 254;
        weight_mem[16'h007F] <= 7;
        weight_mem[16'h0080] <= 242;
        weight_mem[16'h0081] <= 226;
        weight_mem[16'h0082] <= 238;
        weight_mem[16'h0083] <= 247;
        weight_mem[16'h0084] <= 0;
        weight_mem[16'h0085] <= 46;
        weight_mem[16'h0086] <= 59;
        weight_mem[16'h0087] <= 41;
        weight_mem[16'h0088] <= 15;
        weight_mem[16'h0089] <= 27;
        weight_mem[16'h008A] <= 14;
        weight_mem[16'h008B] <= 37;
        weight_mem[16'h008C] <= 47;
        weight_mem[16'h008D] <= 43;
        weight_mem[16'h008E] <= 2;
        weight_mem[16'h008F] <= 9;
        weight_mem[16'h0090] <= 250;
        weight_mem[16'h0091] <= 4;
        weight_mem[16'h0092] <= 236;
        weight_mem[16'h0093] <= 240;
        weight_mem[16'h0094] <= 244;
        weight_mem[16'h0095] <= 241;
        weight_mem[16'h0096] <= 243;
        weight_mem[16'h0097] <= 244;
        weight_mem[16'h0098] <= 226;
        weight_mem[16'h0099] <= 209;
        weight_mem[16'h009A] <= 231;
        weight_mem[16'h009B] <= 245;
        weight_mem[16'h009C] <= 13;
        weight_mem[16'h009D] <= 22;
        weight_mem[16'h009E] <= 15;
        weight_mem[16'h009F] <= 247;
        weight_mem[16'h00A0] <= 240;
        weight_mem[16'h00A1] <= 18;
        weight_mem[16'h00A2] <= 31;
        weight_mem[16'h00A3] <= 47;
        weight_mem[16'h00A4] <= 68;
        weight_mem[16'h00A5] <= 51;
        weight_mem[16'h00A6] <= 13;
        weight_mem[16'h00A7] <= 2;
        weight_mem[16'h00A8] <= 249;
        weight_mem[16'h00A9] <= 251;
        weight_mem[16'h00AA] <= 245;
        weight_mem[16'h00AB] <= 237;
        weight_mem[16'h00AC] <= 251;
        weight_mem[16'h00AD] <= 9;
        weight_mem[16'h00AE] <= 254;
        weight_mem[16'h00AF] <= 240;
        weight_mem[16'h00B0] <= 243;
        weight_mem[16'h00B1] <= 226;
        weight_mem[16'h00B2] <= 4;
        weight_mem[16'h00B3] <= 77;
        weight_mem[16'h00B4] <= 79;
        weight_mem[16'h00B5] <= 15;
        weight_mem[16'h00B6] <= 212;
        weight_mem[16'h00B7] <= 197;
        weight_mem[16'h00B8] <= 225;
        weight_mem[16'h00B9] <= 239;
        weight_mem[16'h00BA] <= 11;
        weight_mem[16'h00BB] <= 13;
        weight_mem[16'h00BC] <= 28;
        weight_mem[16'h00BD] <= 21;
        weight_mem[16'h00BE] <= 14;
        weight_mem[16'h00BF] <= 254;
        weight_mem[16'h00C0] <= 244;
        weight_mem[16'h00C1] <= 254;
        weight_mem[16'h00C2] <= 250;
        weight_mem[16'h00C3] <= 233;
        weight_mem[16'h00C4] <= 255;
        weight_mem[16'h00C5] <= 12;
        weight_mem[16'h00C6] <= 252;
        weight_mem[16'h00C7] <= 2;
        weight_mem[16'h00C8] <= 5;
        weight_mem[16'h00C9] <= 241;
        weight_mem[16'h00CA] <= 34;
        weight_mem[16'h00CB] <= 99;
        weight_mem[16'h00CC] <= 59;
        weight_mem[16'h00CD] <= 212;
        weight_mem[16'h00CE] <= 178;
        weight_mem[16'h00CF] <= 195;
        weight_mem[16'h00D0] <= 214;
        weight_mem[16'h00D1] <= 216;
        weight_mem[16'h00D2] <= 221;
        weight_mem[16'h00D3] <= 244;
        weight_mem[16'h00D4] <= 253;
        weight_mem[16'h00D5] <= 252;
        weight_mem[16'h00D6] <= 8;
        weight_mem[16'h00D7] <= 244;
        weight_mem[16'h00D8] <= 250;
        weight_mem[16'h00D9] <= 2;
        weight_mem[16'h00DA] <= 3;
        weight_mem[16'h00DB] <= 241;
        weight_mem[16'h00DC] <= 253;
        weight_mem[16'h00DD] <= 10;
        weight_mem[16'h00DE] <= 7;
        weight_mem[16'h00DF] <= 253;
        weight_mem[16'h00E0] <= 12;
        weight_mem[16'h00E1] <= 19;
        weight_mem[16'h00E2] <= 71;
        weight_mem[16'h00E3] <= 83;
        weight_mem[16'h00E4] <= 18;
        weight_mem[16'h00E5] <= 185;
        weight_mem[16'h00E6] <= 158;
        weight_mem[16'h00E7] <= 179;
        weight_mem[16'h00E8] <= 197;
        weight_mem[16'h00E9] <= 206;
        weight_mem[16'h00EA] <= 219;
        weight_mem[16'h00EB] <= 224;
        weight_mem[16'h00EC] <= 250;
        weight_mem[16'h00ED] <= 239;
        weight_mem[16'h00EE] <= 242;
        weight_mem[16'h00EF] <= 247;
        weight_mem[16'h00F0] <= 251;
        weight_mem[16'h00F1] <= 2;
        weight_mem[16'h00F2] <= 252;
        weight_mem[16'h00F3] <= 253;
        weight_mem[16'h00F4] <= 6;
        weight_mem[16'h00F5] <= 237;
        weight_mem[16'h00F6] <= 224;
        weight_mem[16'h00F7] <= 253;
        weight_mem[16'h00F8] <= 30;
        weight_mem[16'h00F9] <= 48;
        weight_mem[16'h00FA] <= 81;
        weight_mem[16'h00FB] <= 40;
        weight_mem[16'h00FC] <= 197;
        weight_mem[16'h00FD] <= 144;
        weight_mem[16'h00FE] <= 129;
        weight_mem[16'h00FF] <= 182;
        weight_mem[16'h0100] <= 202;
        weight_mem[16'h0101] <= 209;
        weight_mem[16'h0102] <= 216;
        weight_mem[16'h0103] <= 235;
        weight_mem[16'h0104] <= 249;
        weight_mem[16'h0105] <= 246;
        weight_mem[16'h0106] <= 246;
        weight_mem[16'h0107] <= 242;
        weight_mem[16'h0108] <= 6;
        weight_mem[16'h0109] <= 247;
        weight_mem[16'h010A] <= 253;
        weight_mem[16'h010B] <= 255;
        weight_mem[16'h010C] <= 9;
        weight_mem[16'h010D] <= 251;
        weight_mem[16'h010E] <= 250;
        weight_mem[16'h010F] <= 12;
        weight_mem[16'h0110] <= 54;
        weight_mem[16'h0111] <= 45;
        weight_mem[16'h0112] <= 24;
        weight_mem[16'h0113] <= 217;
        weight_mem[16'h0114] <= 152;
        weight_mem[16'h0115] <= 171;
        weight_mem[16'h0116] <= 190;
        weight_mem[16'h0117] <= 222;
        weight_mem[16'h0118] <= 246;
        weight_mem[16'h0119] <= 250;
        weight_mem[16'h011A] <= 244;
        weight_mem[16'h011B] <= 243;
        weight_mem[16'h011C] <= 240;
        weight_mem[16'h011D] <= 230;
        weight_mem[16'h011E] <= 254;
        weight_mem[16'h011F] <= 3;
        weight_mem[16'h0120] <= 5;
        weight_mem[16'h0121] <= 249;
        weight_mem[16'h0122] <= 255;
        weight_mem[16'h0123] <= 13;
        weight_mem[16'h0124] <= 15;
        weight_mem[16'h0125] <= 40;
        weight_mem[16'h0126] <= 48;
        weight_mem[16'h0127] <= 72;
        weight_mem[16'h0128] <= 82;
        weight_mem[16'h0129] <= 44;
        weight_mem[16'h012A] <= 9;
        weight_mem[16'h012B] <= 225;
        weight_mem[16'h012C] <= 186;
        weight_mem[16'h012D] <= 199;
        weight_mem[16'h012E] <= 244;
        weight_mem[16'h012F] <= 17;
        weight_mem[16'h0130] <= 18;
        weight_mem[16'h0131] <= 20;
        weight_mem[16'h0132] <= 26;
        weight_mem[16'h0133] <= 17;
        weight_mem[16'h0134] <= 1;
        weight_mem[16'h0135] <= 254;
        weight_mem[16'h0136] <= 241;
        weight_mem[16'h0137] <= 249;
        weight_mem[16'h0138] <= 242;
        weight_mem[16'h0139] <= 250;
        weight_mem[16'h013A] <= 3;
        weight_mem[16'h013B] <= 13;
        weight_mem[16'h013C] <= 19;
        weight_mem[16'h013D] <= 57;
        weight_mem[16'h013E] <= 51;
        weight_mem[16'h013F] <= 58;
        weight_mem[16'h0140] <= 55;
        weight_mem[16'h0141] <= 41;
        weight_mem[16'h0142] <= 23;
        weight_mem[16'h0143] <= 0;
        weight_mem[16'h0144] <= 228;
        weight_mem[16'h0145] <= 2;
        weight_mem[16'h0146] <= 16;
        weight_mem[16'h0147] <= 43;
        weight_mem[16'h0148] <= 51;
        weight_mem[16'h0149] <= 39;
        weight_mem[16'h014A] <= 28;
        weight_mem[16'h014B] <= 16;
        weight_mem[16'h014C] <= 8;
        weight_mem[16'h014D] <= 238;
        weight_mem[16'h014E] <= 252;
        weight_mem[16'h014F] <= 253;
        weight_mem[16'h0150] <= 245;
        weight_mem[16'h0151] <= 247;
        weight_mem[16'h0152] <= 4;
        weight_mem[16'h0153] <= 16;
        weight_mem[16'h0154] <= 18;
        weight_mem[16'h0155] <= 22;
        weight_mem[16'h0156] <= 7;
        weight_mem[16'h0157] <= 16;
        weight_mem[16'h0158] <= 14;
        weight_mem[16'h0159] <= 23;
        weight_mem[16'h015A] <= 32;
        weight_mem[16'h015B] <= 41;
        weight_mem[16'h015C] <= 48;
        weight_mem[16'h015D] <= 38;
        weight_mem[16'h015E] <= 60;
        weight_mem[16'h015F] <= 49;
        weight_mem[16'h0160] <= 48;
        weight_mem[16'h0161] <= 22;
        weight_mem[16'h0162] <= 24;
        weight_mem[16'h0163] <= 22;
        weight_mem[16'h0164] <= 254;
        weight_mem[16'h0165] <= 246;
        weight_mem[16'h0166] <= 249;
        weight_mem[16'h0167] <= 6;
        weight_mem[16'h0168] <= 255;
        weight_mem[16'h0169] <= 250;
        weight_mem[16'h016A] <= 245;
        weight_mem[16'h016B] <= 252;
        weight_mem[16'h016C] <= 11;
        weight_mem[16'h016D] <= 253;
        weight_mem[16'h016E] <= 241;
        weight_mem[16'h016F] <= 1;
        weight_mem[16'h0170] <= 17;
        weight_mem[16'h0171] <= 19;
        weight_mem[16'h0172] <= 25;
        weight_mem[16'h0173] <= 38;
        weight_mem[16'h0174] <= 46;
        weight_mem[16'h0175] <= 40;
        weight_mem[16'h0176] <= 47;
        weight_mem[16'h0177] <= 23;
        weight_mem[16'h0178] <= 24;
        weight_mem[16'h0179] <= 24;
        weight_mem[16'h017A] <= 0;
        weight_mem[16'h017B] <= 6;
        weight_mem[16'h017C] <= 249;
        weight_mem[16'h017D] <= 251;
        weight_mem[16'h017E] <= 242;
        weight_mem[16'h017F] <= 252;
        weight_mem[16'h0180] <= 6;
        weight_mem[16'h0181] <= 5;
        weight_mem[16'h0182] <= 6;
        weight_mem[16'h0183] <= 246;
        weight_mem[16'h0184] <= 239;
        weight_mem[16'h0185] <= 234;
        weight_mem[16'h0186] <= 245;
        weight_mem[16'h0187] <= 243;
        weight_mem[16'h0188] <= 244;
        weight_mem[16'h0189] <= 251;
        weight_mem[16'h018A] <= 240;
        weight_mem[16'h018B] <= 3;
        weight_mem[16'h018C] <= 245;
        weight_mem[16'h018D] <= 3;
        weight_mem[16'h018E] <= 3;
        weight_mem[16'h018F] <= 15;
        weight_mem[16'h0190] <= 9;
        weight_mem[16'h0191] <= 3;
        weight_mem[16'h0192] <= 7;
        weight_mem[16'h0193] <= 12;
        weight_mem[16'h0194] <= 249;
        weight_mem[16'h0195] <= 242;
        weight_mem[16'h0196] <= 254;
        weight_mem[16'h0197] <= 242;
        weight_mem[16'h0198] <= 245;
        weight_mem[16'h0199] <= 240;
        weight_mem[16'h019A] <= 244;
        weight_mem[16'h019B] <= 2;
        weight_mem[16'h019C] <= 240;
        weight_mem[16'h019D] <= 3;
        weight_mem[16'h019E] <= 241;
        weight_mem[16'h019F] <= 247;
        weight_mem[16'h01A0] <= 238;
        weight_mem[16'h01A1] <= 250;
        weight_mem[16'h01A2] <= 242;
        weight_mem[16'h01A3] <= 237;
        weight_mem[16'h01A4] <= 248;
        weight_mem[16'h01A5] <= 242;
        weight_mem[16'h01A6] <= 240;
        weight_mem[16'h01A7] <= 1;
        weight_mem[16'h01A8] <= 1;
        weight_mem[16'h01A9] <= 247;
        weight_mem[16'h01AA] <= 253;
        weight_mem[16'h01AB] <= 243;
        weight_mem[16'h01AC] <= 1;
        weight_mem[16'h01AD] <= 251;
        weight_mem[16'h01AE] <= 250;
        weight_mem[16'h01AF] <= 7;

        // layer 1 neuron 1
        weight_mem[16'h0200] <= 0;
        weight_mem[16'h0201] <= 0;
        weight_mem[16'h0202] <= 0;
        weight_mem[16'h0203] <= 0;
        weight_mem[16'h0204] <= 0;
        weight_mem[16'h0205] <= 0;
        weight_mem[16'h0206] <= 0;
        weight_mem[16'h0207] <= 0;
        weight_mem[16'h0208] <= 0;
        weight_mem[16'h0209] <= 0;
        weight_mem[16'h020A] <= 0;
        weight_mem[16'h020B] <= 0;
        weight_mem[16'h020C] <= 0;
        weight_mem[16'h020D] <= 0;
        weight_mem[16'h020E] <= 0;
        weight_mem[16'h020F] <= 0;
        weight_mem[16'h0210] <= 0;
        weight_mem[16'h0211] <= 0;
        weight_mem[16'h0212] <= 0;
        weight_mem[16'h0213] <= 0;
        weight_mem[16'h0214] <= 0;
        weight_mem[16'h0215] <= 0;
        weight_mem[16'h0216] <= 0;
        weight_mem[16'h0217] <= 0;
        weight_mem[16'h0218] <= 0;
        weight_mem[16'h0219] <= 0;
        weight_mem[16'h021A] <= 0;
        weight_mem[16'h021B] <= 0;
        weight_mem[16'h021C] <= 0;
        weight_mem[16'h021D] <= 0;
        weight_mem[16'h021E] <= 0;
        weight_mem[16'h021F] <= 0;
        weight_mem[16'h0220] <= 0;
        weight_mem[16'h0221] <= 0;
        weight_mem[16'h0222] <= 0;
        weight_mem[16'h0223] <= 0;
        weight_mem[16'h0224] <= 0;
        weight_mem[16'h0225] <= 0;
        weight_mem[16'h0226] <= 0;
        weight_mem[16'h0227] <= 0;
        weight_mem[16'h0228] <= 0;
        weight_mem[16'h0229] <= 0;
        weight_mem[16'h022A] <= 0;
        weight_mem[16'h022B] <= 0;
        weight_mem[16'h022C] <= 0;
        weight_mem[16'h022D] <= 0;
        weight_mem[16'h022E] <= 0;
        weight_mem[16'h022F] <= 0;
        weight_mem[16'h0230] <= 0;
        weight_mem[16'h0231] <= 0;
        weight_mem[16'h0232] <= 0;
        weight_mem[16'h0233] <= 0;
        weight_mem[16'h0234] <= 0;
        weight_mem[16'h0235] <= 0;
        weight_mem[16'h0236] <= 0;
        weight_mem[16'h0237] <= 0;
        weight_mem[16'h0238] <= 0;
        weight_mem[16'h0239] <= 0;
        weight_mem[16'h023A] <= 0;
        weight_mem[16'h023B] <= 0;
        weight_mem[16'h023C] <= 0;
        weight_mem[16'h023D] <= 0;
        weight_mem[16'h023E] <= 0;
        weight_mem[16'h023F] <= 0;
        weight_mem[16'h0240] <= 0;
        weight_mem[16'h0241] <= 0;
        weight_mem[16'h0242] <= 0;
        weight_mem[16'h0243] <= 0;
        weight_mem[16'h0244] <= 0;
        weight_mem[16'h0245] <= 0;
        weight_mem[16'h0246] <= 0;
        weight_mem[16'h0247] <= 0;
        weight_mem[16'h0248] <= 0;
        weight_mem[16'h0249] <= 0;
        weight_mem[16'h024A] <= 0;
        weight_mem[16'h024B] <= 0;
        weight_mem[16'h024C] <= 0;
        weight_mem[16'h024D] <= 0;
        weight_mem[16'h024E] <= 0;
        weight_mem[16'h024F] <= 0;
        weight_mem[16'h0250] <= 0;
        weight_mem[16'h0251] <= 0;
        weight_mem[16'h0252] <= 0;
        weight_mem[16'h0253] <= 0;
        weight_mem[16'h0254] <= 0;
        weight_mem[16'h0255] <= 0;
        weight_mem[16'h0256] <= 0;
        weight_mem[16'h0257] <= 0;
        weight_mem[16'h0258] <= 0;
        weight_mem[16'h0259] <= 0;
        weight_mem[16'h025A] <= 0;
        weight_mem[16'h025B] <= 0;
        weight_mem[16'h025C] <= 0;
        weight_mem[16'h025D] <= 0;
        weight_mem[16'h025E] <= 0;
        weight_mem[16'h025F] <= 0;
        weight_mem[16'h0260] <= 0;
        weight_mem[16'h0261] <= 0;
        weight_mem[16'h0262] <= 0;
        weight_mem[16'h0263] <= 0;
        weight_mem[16'h0264] <= 0;
        weight_mem[16'h0265] <= 0;
        weight_mem[16'h0266] <= 0;
        weight_mem[16'h0267] <= 0;
        weight_mem[16'h0268] <= 0;
        weight_mem[16'h0269] <= 0;
        weight_mem[16'h026A] <= 0;
        weight_mem[16'h026B] <= 0;
        weight_mem[16'h026C] <= 0;
        weight_mem[16'h026D] <= 0;
        weight_mem[16'h026E] <= 0;
        weight_mem[16'h026F] <= 0;
        weight_mem[16'h0270] <= 0;
        weight_mem[16'h0271] <= 0;
        weight_mem[16'h0272] <= 0;
        weight_mem[16'h0273] <= 0;
        weight_mem[16'h0274] <= 0;
        weight_mem[16'h0275] <= 0;
        weight_mem[16'h0276] <= 0;
        weight_mem[16'h0277] <= 0;
        weight_mem[16'h0278] <= 0;
        weight_mem[16'h0279] <= 0;
        weight_mem[16'h027A] <= 0;
        weight_mem[16'h027B] <= 0;
        weight_mem[16'h027C] <= 0;
        weight_mem[16'h027D] <= 0;
        weight_mem[16'h027E] <= 0;
        weight_mem[16'h027F] <= 0;
        weight_mem[16'h0280] <= 0;
        weight_mem[16'h0281] <= 0;
        weight_mem[16'h0282] <= 0;
        weight_mem[16'h0283] <= 0;
        weight_mem[16'h0284] <= 0;
        weight_mem[16'h0285] <= 0;
        weight_mem[16'h0286] <= 0;
        weight_mem[16'h0287] <= 0;
        weight_mem[16'h0288] <= 0;
        weight_mem[16'h0289] <= 0;
        weight_mem[16'h028A] <= 0;
        weight_mem[16'h028B] <= 0;
        weight_mem[16'h028C] <= 0;
        weight_mem[16'h028D] <= 0;
        weight_mem[16'h028E] <= 0;
        weight_mem[16'h028F] <= 0;
        weight_mem[16'h0290] <= 0;
        weight_mem[16'h0291] <= 0;
        weight_mem[16'h0292] <= 0;
        weight_mem[16'h0293] <= 0;
        weight_mem[16'h0294] <= 0;
        weight_mem[16'h0295] <= 0;
        weight_mem[16'h0296] <= 0;
        weight_mem[16'h0297] <= 0;
        weight_mem[16'h0298] <= 0;
        weight_mem[16'h0299] <= 0;
        weight_mem[16'h029A] <= 0;
        weight_mem[16'h029B] <= 0;
        weight_mem[16'h029C] <= 0;
        weight_mem[16'h029D] <= 0;
        weight_mem[16'h029E] <= 0;
        weight_mem[16'h029F] <= 0;
        weight_mem[16'h02A0] <= 0;
        weight_mem[16'h02A1] <= 0;
        weight_mem[16'h02A2] <= 0;
        weight_mem[16'h02A3] <= 0;
        weight_mem[16'h02A4] <= 0;
        weight_mem[16'h02A5] <= 0;
        weight_mem[16'h02A6] <= 0;
        weight_mem[16'h02A7] <= 0;
        weight_mem[16'h02A8] <= 0;
        weight_mem[16'h02A9] <= 0;
        weight_mem[16'h02AA] <= 0;
        weight_mem[16'h02AB] <= 0;
        weight_mem[16'h02AC] <= 0;
        weight_mem[16'h02AD] <= 0;
        weight_mem[16'h02AE] <= 0;
        weight_mem[16'h02AF] <= 0;
        weight_mem[16'h02B0] <= 0;
        weight_mem[16'h02B1] <= 0;
        weight_mem[16'h02B2] <= 0;
        weight_mem[16'h02B3] <= 0;
        weight_mem[16'h02B4] <= 0;
        weight_mem[16'h02B5] <= 0;
        weight_mem[16'h02B6] <= 0;
        weight_mem[16'h02B7] <= 0;
        weight_mem[16'h02B8] <= 0;
        weight_mem[16'h02B9] <= 0;
        weight_mem[16'h02BA] <= 0;
        weight_mem[16'h02BB] <= 0;
        weight_mem[16'h02BC] <= 0;
        weight_mem[16'h02BD] <= 0;
        weight_mem[16'h02BE] <= 0;
        weight_mem[16'h02BF] <= 0;
        weight_mem[16'h02C0] <= 0;
        weight_mem[16'h02C1] <= 0;
        weight_mem[16'h02C2] <= 0;
        weight_mem[16'h02C3] <= 0;
        weight_mem[16'h02C4] <= 0;
        weight_mem[16'h02C5] <= 0;
        weight_mem[16'h02C6] <= 0;
        weight_mem[16'h02C7] <= 0;
        weight_mem[16'h02C8] <= 0;
        weight_mem[16'h02C9] <= 0;
        weight_mem[16'h02CA] <= 0;
        weight_mem[16'h02CB] <= 0;
        weight_mem[16'h02CC] <= 0;
        weight_mem[16'h02CD] <= 0;
        weight_mem[16'h02CE] <= 0;
        weight_mem[16'h02CF] <= 0;
        weight_mem[16'h02D0] <= 0;
        weight_mem[16'h02D1] <= 0;
        weight_mem[16'h02D2] <= 0;
        weight_mem[16'h02D3] <= 0;
        weight_mem[16'h02D4] <= 0;
        weight_mem[16'h02D5] <= 0;
        weight_mem[16'h02D6] <= 0;
        weight_mem[16'h02D7] <= 0;
        weight_mem[16'h02D8] <= 0;
        weight_mem[16'h02D9] <= 0;
        weight_mem[16'h02DA] <= 0;
        weight_mem[16'h02DB] <= 0;
        weight_mem[16'h02DC] <= 0;
        weight_mem[16'h02DD] <= 0;
        weight_mem[16'h02DE] <= 0;
        weight_mem[16'h02DF] <= 0;
        weight_mem[16'h02E0] <= 0;
        weight_mem[16'h02E1] <= 0;
        weight_mem[16'h02E2] <= 0;
        weight_mem[16'h02E3] <= 255;
        weight_mem[16'h02E4] <= 255;
        weight_mem[16'h02E5] <= 0;
        weight_mem[16'h02E6] <= 0;
        weight_mem[16'h02E7] <= 0;
        weight_mem[16'h02E8] <= 0;
        weight_mem[16'h02E9] <= 0;
        weight_mem[16'h02EA] <= 0;
        weight_mem[16'h02EB] <= 0;
        weight_mem[16'h02EC] <= 0;
        weight_mem[16'h02ED] <= 0;
        weight_mem[16'h02EE] <= 0;
        weight_mem[16'h02EF] <= 0;
        weight_mem[16'h02F0] <= 0;
        weight_mem[16'h02F1] <= 0;
        weight_mem[16'h02F2] <= 0;
        weight_mem[16'h02F3] <= 0;
        weight_mem[16'h02F4] <= 0;
        weight_mem[16'h02F5] <= 0;
        weight_mem[16'h02F6] <= 0;
        weight_mem[16'h02F7] <= 0;
        weight_mem[16'h02F8] <= 0;
        weight_mem[16'h02F9] <= 0;
        weight_mem[16'h02FA] <= 0;
        weight_mem[16'h02FB] <= 255;
        weight_mem[16'h02FC] <= 0;
        weight_mem[16'h02FD] <= 0;
        weight_mem[16'h02FE] <= 0;
        weight_mem[16'h02FF] <= 0;
        weight_mem[16'h0300] <= 0;
        weight_mem[16'h0301] <= 0;
        weight_mem[16'h0302] <= 0;
        weight_mem[16'h0303] <= 0;
        weight_mem[16'h0304] <= 0;
        weight_mem[16'h0305] <= 0;
        weight_mem[16'h0306] <= 0;
        weight_mem[16'h0307] <= 0;
        weight_mem[16'h0308] <= 0;
        weight_mem[16'h0309] <= 0;
        weight_mem[16'h030A] <= 0;
        weight_mem[16'h030B] <= 0;
        weight_mem[16'h030C] <= 0;
        weight_mem[16'h030D] <= 0;
        weight_mem[16'h030E] <= 0;
        weight_mem[16'h030F] <= 0;
        weight_mem[16'h0310] <= 0;
        weight_mem[16'h0311] <= 0;
        weight_mem[16'h0312] <= 0;
        weight_mem[16'h0313] <= 0;
        weight_mem[16'h0314] <= 0;
        weight_mem[16'h0315] <= 0;
        weight_mem[16'h0316] <= 0;
        weight_mem[16'h0317] <= 0;
        weight_mem[16'h0318] <= 0;
        weight_mem[16'h0319] <= 0;
        weight_mem[16'h031A] <= 0;
        weight_mem[16'h031B] <= 0;
        weight_mem[16'h031C] <= 0;
        weight_mem[16'h031D] <= 0;
        weight_mem[16'h031E] <= 0;
        weight_mem[16'h031F] <= 0;
        weight_mem[16'h0320] <= 0;
        weight_mem[16'h0321] <= 0;
        weight_mem[16'h0322] <= 0;
        weight_mem[16'h0323] <= 0;
        weight_mem[16'h0324] <= 0;
        weight_mem[16'h0325] <= 0;
        weight_mem[16'h0326] <= 0;
        weight_mem[16'h0327] <= 0;
        weight_mem[16'h0328] <= 0;
        weight_mem[16'h0329] <= 0;
        weight_mem[16'h032A] <= 0;
        weight_mem[16'h032B] <= 0;
        weight_mem[16'h032C] <= 0;
        weight_mem[16'h032D] <= 0;
        weight_mem[16'h032E] <= 0;
        weight_mem[16'h032F] <= 0;
        weight_mem[16'h0330] <= 0;
        weight_mem[16'h0331] <= 0;
        weight_mem[16'h0332] <= 0;
        weight_mem[16'h0333] <= 0;
        weight_mem[16'h0334] <= 0;
        weight_mem[16'h0335] <= 0;
        weight_mem[16'h0336] <= 0;
        weight_mem[16'h0337] <= 0;
        weight_mem[16'h0338] <= 0;
        weight_mem[16'h0339] <= 0;
        weight_mem[16'h033A] <= 0;
        weight_mem[16'h033B] <= 0;
        weight_mem[16'h033C] <= 0;
        weight_mem[16'h033D] <= 0;
        weight_mem[16'h033E] <= 0;
        weight_mem[16'h033F] <= 0;
        weight_mem[16'h0340] <= 0;
        weight_mem[16'h0341] <= 0;
        weight_mem[16'h0342] <= 0;
        weight_mem[16'h0343] <= 0;
        weight_mem[16'h0344] <= 0;
        weight_mem[16'h0345] <= 0;
        weight_mem[16'h0346] <= 0;
        weight_mem[16'h0347] <= 0;
        weight_mem[16'h0348] <= 0;
        weight_mem[16'h0349] <= 0;
        weight_mem[16'h034A] <= 0;
        weight_mem[16'h034B] <= 0;
        weight_mem[16'h034C] <= 0;
        weight_mem[16'h034D] <= 0;
        weight_mem[16'h034E] <= 0;
        weight_mem[16'h034F] <= 0;
        weight_mem[16'h0350] <= 0;
        weight_mem[16'h0351] <= 0;
        weight_mem[16'h0352] <= 0;
        weight_mem[16'h0353] <= 0;
        weight_mem[16'h0354] <= 0;
        weight_mem[16'h0355] <= 0;
        weight_mem[16'h0356] <= 0;
        weight_mem[16'h0357] <= 0;
        weight_mem[16'h0358] <= 0;
        weight_mem[16'h0359] <= 0;
        weight_mem[16'h035A] <= 0;
        weight_mem[16'h035B] <= 0;
        weight_mem[16'h035C] <= 0;
        weight_mem[16'h035D] <= 0;
        weight_mem[16'h035E] <= 0;
        weight_mem[16'h035F] <= 0;
        weight_mem[16'h0360] <= 0;
        weight_mem[16'h0361] <= 0;
        weight_mem[16'h0362] <= 0;
        weight_mem[16'h0363] <= 0;
        weight_mem[16'h0364] <= 0;
        weight_mem[16'h0365] <= 0;
        weight_mem[16'h0366] <= 0;
        weight_mem[16'h0367] <= 0;
        weight_mem[16'h0368] <= 0;
        weight_mem[16'h0369] <= 0;
        weight_mem[16'h036A] <= 0;
        weight_mem[16'h036B] <= 0;
        weight_mem[16'h036C] <= 0;
        weight_mem[16'h036D] <= 0;
        weight_mem[16'h036E] <= 0;
        weight_mem[16'h036F] <= 0;
        weight_mem[16'h0370] <= 0;
        weight_mem[16'h0371] <= 0;
        weight_mem[16'h0372] <= 0;
        weight_mem[16'h0373] <= 0;
        weight_mem[16'h0374] <= 0;
        weight_mem[16'h0375] <= 0;
        weight_mem[16'h0376] <= 0;
        weight_mem[16'h0377] <= 0;
        weight_mem[16'h0378] <= 0;
        weight_mem[16'h0379] <= 0;
        weight_mem[16'h037A] <= 0;
        weight_mem[16'h037B] <= 0;
        weight_mem[16'h037C] <= 0;
        weight_mem[16'h037D] <= 0;
        weight_mem[16'h037E] <= 0;
        weight_mem[16'h037F] <= 0;
        weight_mem[16'h0380] <= 0;
        weight_mem[16'h0381] <= 0;
        weight_mem[16'h0382] <= 0;
        weight_mem[16'h0383] <= 0;
        weight_mem[16'h0384] <= 0;
        weight_mem[16'h0385] <= 0;
        weight_mem[16'h0386] <= 0;
        weight_mem[16'h0387] <= 0;
        weight_mem[16'h0388] <= 0;
        weight_mem[16'h0389] <= 0;
        weight_mem[16'h038A] <= 0;
        weight_mem[16'h038B] <= 0;
        weight_mem[16'h038C] <= 0;
        weight_mem[16'h038D] <= 0;
        weight_mem[16'h038E] <= 0;
        weight_mem[16'h038F] <= 0;
        weight_mem[16'h0390] <= 0;
        weight_mem[16'h0391] <= 0;
        weight_mem[16'h0392] <= 0;
        weight_mem[16'h0393] <= 0;
        weight_mem[16'h0394] <= 0;
        weight_mem[16'h0395] <= 0;
        weight_mem[16'h0396] <= 0;
        weight_mem[16'h0397] <= 0;
        weight_mem[16'h0398] <= 0;
        weight_mem[16'h0399] <= 0;
        weight_mem[16'h039A] <= 0;
        weight_mem[16'h039B] <= 0;
        weight_mem[16'h039C] <= 0;
        weight_mem[16'h039D] <= 0;
        weight_mem[16'h039E] <= 0;
        weight_mem[16'h039F] <= 0;
        weight_mem[16'h03A0] <= 0;
        weight_mem[16'h03A1] <= 0;
        weight_mem[16'h03A2] <= 0;
        weight_mem[16'h03A3] <= 0;
        weight_mem[16'h03A4] <= 0;
        weight_mem[16'h03A5] <= 0;
        weight_mem[16'h03A6] <= 0;
        weight_mem[16'h03A7] <= 0;
        weight_mem[16'h03A8] <= 0;
        weight_mem[16'h03A9] <= 0;
        weight_mem[16'h03AA] <= 0;
        weight_mem[16'h03AB] <= 0;
        weight_mem[16'h03AC] <= 0;
        weight_mem[16'h03AD] <= 0;
        weight_mem[16'h03AE] <= 0;
        weight_mem[16'h03AF] <= 0;

        // layer 1 neuron 2
        weight_mem[16'h0400] <= 179;
        weight_mem[16'h0401] <= 179;
        weight_mem[16'h0402] <= 179;
        weight_mem[16'h0403] <= 179;
        weight_mem[16'h0404] <= 179;
        weight_mem[16'h0405] <= 179;
        weight_mem[16'h0406] <= 179;
        weight_mem[16'h0407] <= 179;
        weight_mem[16'h0408] <= 179;
        weight_mem[16'h0409] <= 179;
        weight_mem[16'h040A] <= 179;
        weight_mem[16'h040B] <= 179;
        weight_mem[16'h040C] <= 179;
        weight_mem[16'h040D] <= 179;
        weight_mem[16'h040E] <= 179;
        weight_mem[16'h040F] <= 179;
        weight_mem[16'h0410] <= 179;
        weight_mem[16'h0411] <= 179;
        weight_mem[16'h0412] <= 179;
        weight_mem[16'h0413] <= 179;
        weight_mem[16'h0414] <= 179;
        weight_mem[16'h0415] <= 179;
        weight_mem[16'h0416] <= 179;
        weight_mem[16'h0417] <= 179;
        weight_mem[16'h0418] <= 179;
        weight_mem[16'h0419] <= 179;
        weight_mem[16'h041A] <= 179;
        weight_mem[16'h041B] <= 179;
        weight_mem[16'h041C] <= 179;
        weight_mem[16'h041D] <= 179;
        weight_mem[16'h041E] <= 179;
        weight_mem[16'h041F] <= 180;
        weight_mem[16'h0420] <= 180;
        weight_mem[16'h0421] <= 181;
        weight_mem[16'h0422] <= 181;
        weight_mem[16'h0423] <= 179;
        weight_mem[16'h0424] <= 178;
        weight_mem[16'h0425] <= 180;
        weight_mem[16'h0426] <= 182;
        weight_mem[16'h0427] <= 182;
        weight_mem[16'h0428] <= 180;
        weight_mem[16'h0429] <= 181;
        weight_mem[16'h042A] <= 180;
        weight_mem[16'h042B] <= 179;
        weight_mem[16'h042C] <= 179;
        weight_mem[16'h042D] <= 179;
        weight_mem[16'h042E] <= 179;
        weight_mem[16'h042F] <= 179;
        weight_mem[16'h0430] <= 179;
        weight_mem[16'h0431] <= 179;
        weight_mem[16'h0432] <= 179;
        weight_mem[16'h0433] <= 179;
        weight_mem[16'h0434] <= 179;
        weight_mem[16'h0435] <= 180;
        weight_mem[16'h0436] <= 181;
        weight_mem[16'h0437] <= 187;
        weight_mem[16'h0438] <= 196;
        weight_mem[16'h0439] <= 199;
        weight_mem[16'h043A] <= 193;
        weight_mem[16'h043B] <= 188;
        weight_mem[16'h043C] <= 188;
        weight_mem[16'h043D] <= 190;
        weight_mem[16'h043E] <= 199;
        weight_mem[16'h043F] <= 200;
        weight_mem[16'h0440] <= 189;
        weight_mem[16'h0441] <= 187;
        weight_mem[16'h0442] <= 182;
        weight_mem[16'h0443] <= 178;
        weight_mem[16'h0444] <= 179;
        weight_mem[16'h0445] <= 179;
        weight_mem[16'h0446] <= 179;
        weight_mem[16'h0447] <= 179;
        weight_mem[16'h0448] <= 179;
        weight_mem[16'h0449] <= 179;
        weight_mem[16'h044A] <= 179;
        weight_mem[16'h044B] <= 180;
        weight_mem[16'h044C] <= 180;
        weight_mem[16'h044D] <= 179;
        weight_mem[16'h044E] <= 178;
        weight_mem[16'h044F] <= 184;
        weight_mem[16'h0450] <= 194;
        weight_mem[16'h0451] <= 207;
        weight_mem[16'h0452] <= 212;
        weight_mem[16'h0453] <= 197;
        weight_mem[16'h0454] <= 191;
        weight_mem[16'h0455] <= 189;
        weight_mem[16'h0456] <= 189;
        weight_mem[16'h0457] <= 200;
        weight_mem[16'h0458] <= 209;
        weight_mem[16'h0459] <= 210;
        weight_mem[16'h045A] <= 199;
        weight_mem[16'h045B] <= 185;
        weight_mem[16'h045C] <= 175;
        weight_mem[16'h045D] <= 176;
        weight_mem[16'h045E] <= 180;
        weight_mem[16'h045F] <= 180;
        weight_mem[16'h0460] <= 179;
        weight_mem[16'h0461] <= 179;
        weight_mem[16'h0462] <= 179;
        weight_mem[16'h0463] <= 180;
        weight_mem[16'h0464] <= 179;
        weight_mem[16'h0465] <= 174;
        weight_mem[16'h0466] <= 175;
        weight_mem[16'h0467] <= 192;
        weight_mem[16'h0468] <= 204;
        weight_mem[16'h0469] <= 207;
        weight_mem[16'h046A] <= 209;
        weight_mem[16'h046B] <= 190;
        weight_mem[16'h046C] <= 188;
        weight_mem[16'h046D] <= 224;
        weight_mem[16'h046E] <= 243;
        weight_mem[16'h046F] <= 242;
        weight_mem[16'h0470] <= 239;
        weight_mem[16'h0471] <= 227;
        weight_mem[16'h0472] <= 211;
        weight_mem[16'h0473] <= 184;
        weight_mem[16'h0474] <= 174;
        weight_mem[16'h0475] <= 179;
        weight_mem[16'h0476] <= 181;
        weight_mem[16'h0477] <= 180;
        weight_mem[16'h0478] <= 179;
        weight_mem[16'h0479] <= 179;
        weight_mem[16'h047A] <= 178;
        weight_mem[16'h047B] <= 177;
        weight_mem[16'h047C] <= 174;
        weight_mem[16'h047D] <= 173;
        weight_mem[16'h047E] <= 182;
        weight_mem[16'h047F] <= 203;
        weight_mem[16'h0480] <= 215;
        weight_mem[16'h0481] <= 217;
        weight_mem[16'h0482] <= 229;
        weight_mem[16'h0483] <= 227;
        weight_mem[16'h0484] <= 235;
        weight_mem[16'h0485] <= 241;
        weight_mem[16'h0486] <= 1;
        weight_mem[16'h0487] <= 249;
        weight_mem[16'h0488] <= 239;
        weight_mem[16'h0489] <= 232;
        weight_mem[16'h048A] <= 222;
        weight_mem[16'h048B] <= 195;
        weight_mem[16'h048C] <= 189;
        weight_mem[16'h048D] <= 187;
        weight_mem[16'h048E] <= 181;
        weight_mem[16'h048F] <= 180;
        weight_mem[16'h0490] <= 179;
        weight_mem[16'h0491] <= 179;
        weight_mem[16'h0492] <= 178;
        weight_mem[16'h0493] <= 177;
        weight_mem[16'h0494] <= 177;
        weight_mem[16'h0495] <= 189;
        weight_mem[16'h0496] <= 194;
        weight_mem[16'h0497] <= 208;
        weight_mem[16'h0498] <= 226;
        weight_mem[16'h0499] <= 13;
        weight_mem[16'h049A] <= 28;
        weight_mem[16'h049B] <= 17;
        weight_mem[16'h049C] <= 240;
        weight_mem[16'h049D] <= 186;
        weight_mem[16'h049E] <= 182;
        weight_mem[16'h049F] <= 211;
        weight_mem[16'h04A0] <= 216;
        weight_mem[16'h04A1] <= 211;
        weight_mem[16'h04A2] <= 208;
        weight_mem[16'h04A3] <= 212;
        weight_mem[16'h04A4] <= 203;
        weight_mem[16'h04A5] <= 188;
        weight_mem[16'h04A6] <= 180;
        weight_mem[16'h04A7] <= 179;
        weight_mem[16'h04A8] <= 179;
        weight_mem[16'h04A9] <= 179;
        weight_mem[16'h04AA] <= 179;
        weight_mem[16'h04AB] <= 181;
        weight_mem[16'h04AC] <= 190;
        weight_mem[16'h04AD] <= 196;
        weight_mem[16'h04AE] <= 178;
        weight_mem[16'h04AF] <= 163;
        weight_mem[16'h04B0] <= 213;
        weight_mem[16'h04B1] <= 25;
        weight_mem[16'h04B2] <= 29;
        weight_mem[16'h04B3] <= 248;
        weight_mem[16'h04B4] <= 203;
        weight_mem[16'h04B5] <= 162;
        weight_mem[16'h04B6] <= 194;
        weight_mem[16'h04B7] <= 222;
        weight_mem[16'h04B8] <= 207;
        weight_mem[16'h04B9] <= 184;
        weight_mem[16'h04BA] <= 186;
        weight_mem[16'h04BB] <= 205;
        weight_mem[16'h04BC] <= 199;
        weight_mem[16'h04BD] <= 186;
        weight_mem[16'h04BE] <= 179;
        weight_mem[16'h04BF] <= 179;
        weight_mem[16'h04C0] <= 179;
        weight_mem[16'h04C1] <= 179;
        weight_mem[16'h04C2] <= 179;
        weight_mem[16'h04C3] <= 185;
        weight_mem[16'h04C4] <= 185;
        weight_mem[16'h04C5] <= 171;
        weight_mem[16'h04C6] <= 128;
        weight_mem[16'h04C7] <= 130;
        weight_mem[16'h04C8] <= 199;
        weight_mem[16'h04C9] <= 234;
        weight_mem[16'h04CA] <= 226;
        weight_mem[16'h04CB] <= 205;
        weight_mem[16'h04CC] <= 198;
        weight_mem[16'h04CD] <= 195;
        weight_mem[16'h04CE] <= 217;
        weight_mem[16'h04CF] <= 214;
        weight_mem[16'h04D0] <= 193;
        weight_mem[16'h04D1] <= 187;
        weight_mem[16'h04D2] <= 191;
        weight_mem[16'h04D3] <= 201;
        weight_mem[16'h04D4] <= 192;
        weight_mem[16'h04D5] <= 187;
        weight_mem[16'h04D6] <= 185;
        weight_mem[16'h04D7] <= 180;
        weight_mem[16'h04D8] <= 179;
        weight_mem[16'h04D9] <= 179;
        weight_mem[16'h04DA] <= 179;
        weight_mem[16'h04DB] <= 180;
        weight_mem[16'h04DC] <= 179;
        weight_mem[16'h04DD] <= 171;
        weight_mem[16'h04DE] <= 158;
        weight_mem[16'h04DF] <= 198;
        weight_mem[16'h04E0] <= 249;
        weight_mem[16'h04E1] <= 250;
        weight_mem[16'h04E2] <= 232;
        weight_mem[16'h04E3] <= 216;
        weight_mem[16'h04E4] <= 212;
        weight_mem[16'h04E5] <= 215;
        weight_mem[16'h04E6] <= 245;
        weight_mem[16'h04E7] <= 230;
        weight_mem[16'h04E8] <= 198;
        weight_mem[16'h04E9] <= 199;
        weight_mem[16'h04EA] <= 205;
        weight_mem[16'h04EB] <= 209;
        weight_mem[16'h04EC] <= 195;
        weight_mem[16'h04ED] <= 185;
        weight_mem[16'h04EE] <= 186;
        weight_mem[16'h04EF] <= 181;
        weight_mem[16'h04F0] <= 179;
        weight_mem[16'h04F1] <= 179;
        weight_mem[16'h04F2] <= 180;
        weight_mem[16'h04F3] <= 180;
        weight_mem[16'h04F4] <= 183;
        weight_mem[16'h04F5] <= 186;
        weight_mem[16'h04F6] <= 227;
        weight_mem[16'h04F7] <= 22;
        weight_mem[16'h04F8] <= 35;
        weight_mem[16'h04F9] <= 21;
        weight_mem[16'h04FA] <= 250;
        weight_mem[16'h04FB] <= 220;
        weight_mem[16'h04FC] <= 221;
        weight_mem[16'h04FD] <= 227;
        weight_mem[16'h04FE] <= 238;
        weight_mem[16'h04FF] <= 229;
        weight_mem[16'h0500] <= 218;
        weight_mem[16'h0501] <= 213;
        weight_mem[16'h0502] <= 201;
        weight_mem[16'h0503] <= 197;
        weight_mem[16'h0504] <= 183;
        weight_mem[16'h0505] <= 175;
        weight_mem[16'h0506] <= 180;
        weight_mem[16'h0507] <= 181;
        weight_mem[16'h0508] <= 179;
        weight_mem[16'h0509] <= 179;
        weight_mem[16'h050A] <= 186;
        weight_mem[16'h050B] <= 194;
        weight_mem[16'h050C] <= 199;
        weight_mem[16'h050D] <= 203;
        weight_mem[16'h050E] <= 220;
        weight_mem[16'h050F] <= 242;
        weight_mem[16'h0510] <= 250;
        weight_mem[16'h0511] <= 253;
        weight_mem[16'h0512] <= 253;
        weight_mem[16'h0513] <= 237;
        weight_mem[16'h0514] <= 217;
        weight_mem[16'h0515] <= 211;
        weight_mem[16'h0516] <= 216;
        weight_mem[16'h0517] <= 211;
        weight_mem[16'h0518] <= 218;
        weight_mem[16'h0519] <= 206;
        weight_mem[16'h051A] <= 192;
        weight_mem[16'h051B] <= 185;
        weight_mem[16'h051C] <= 181;
        weight_mem[16'h051D] <= 181;
        weight_mem[16'h051E] <= 183;
        weight_mem[16'h051F] <= 181;
        weight_mem[16'h0520] <= 179;
        weight_mem[16'h0521] <= 179;
        weight_mem[16'h0522] <= 182;
        weight_mem[16'h0523] <= 187;
        weight_mem[16'h0524] <= 194;
        weight_mem[16'h0525] <= 205;
        weight_mem[16'h0526] <= 217;
        weight_mem[16'h0527] <= 234;
        weight_mem[16'h0528] <= 250;
        weight_mem[16'h0529] <= 255;
        weight_mem[16'h052A] <= 249;
        weight_mem[16'h052B] <= 227;
        weight_mem[16'h052C] <= 192;
        weight_mem[16'h052D] <= 183;
        weight_mem[16'h052E] <= 194;
        weight_mem[16'h052F] <= 209;
        weight_mem[16'h0530] <= 234;
        weight_mem[16'h0531] <= 211;
        weight_mem[16'h0532] <= 179;
        weight_mem[16'h0533] <= 176;
        weight_mem[16'h0534] <= 175;
        weight_mem[16'h0535] <= 178;
        weight_mem[16'h0536] <= 179;
        weight_mem[16'h0537] <= 179;
        weight_mem[16'h0538] <= 179;
        weight_mem[16'h0539] <= 179;
        weight_mem[16'h053A] <= 180;
        weight_mem[16'h053B] <= 178;
        weight_mem[16'h053C] <= 164;
        weight_mem[16'h053D] <= 170;
        weight_mem[16'h053E] <= 206;
        weight_mem[16'h053F] <= 236;
        weight_mem[16'h0540] <= 0;
        weight_mem[16'h0541] <= 5;
        weight_mem[16'h0542] <= 1;
        weight_mem[16'h0543] <= 235;
        weight_mem[16'h0544] <= 200;
        weight_mem[16'h0545] <= 216;
        weight_mem[16'h0546] <= 220;
        weight_mem[16'h0547] <= 213;
        weight_mem[16'h0548] <= 223;
        weight_mem[16'h0549] <= 191;
        weight_mem[16'h054A] <= 171;
        weight_mem[16'h054B] <= 175;
        weight_mem[16'h054C] <= 178;
        weight_mem[16'h054D] <= 180;
        weight_mem[16'h054E] <= 180;
        weight_mem[16'h054F] <= 179;
        weight_mem[16'h0550] <= 179;
        weight_mem[16'h0551] <= 179;
        weight_mem[16'h0552] <= 180;
        weight_mem[16'h0553] <= 180;
        weight_mem[16'h0554] <= 168;
        weight_mem[16'h0555] <= 168;
        weight_mem[16'h0556] <= 197;
        weight_mem[16'h0557] <= 223;
        weight_mem[16'h0558] <= 224;
        weight_mem[16'h0559] <= 229;
        weight_mem[16'h055A] <= 228;
        weight_mem[16'h055B] <= 226;
        weight_mem[16'h055C] <= 234;
        weight_mem[16'h055D] <= 233;
        weight_mem[16'h055E] <= 201;
        weight_mem[16'h055F] <= 180;
        weight_mem[16'h0560] <= 183;
        weight_mem[16'h0561] <= 177;
        weight_mem[16'h0562] <= 177;
        weight_mem[16'h0563] <= 179;
        weight_mem[16'h0564] <= 179;
        weight_mem[16'h0565] <= 178;
        weight_mem[16'h0566] <= 179;
        weight_mem[16'h0567] <= 179;
        weight_mem[16'h0568] <= 179;
        weight_mem[16'h0569] <= 179;
        weight_mem[16'h056A] <= 180;
        weight_mem[16'h056B] <= 183;
        weight_mem[16'h056C] <= 182;
        weight_mem[16'h056D] <= 184;
        weight_mem[16'h056E] <= 194;
        weight_mem[16'h056F] <= 200;
        weight_mem[16'h0570] <= 198;
        weight_mem[16'h0571] <= 196;
        weight_mem[16'h0572] <= 195;
        weight_mem[16'h0573] <= 193;
        weight_mem[16'h0574] <= 202;
        weight_mem[16'h0575] <= 195;
        weight_mem[16'h0576] <= 186;
        weight_mem[16'h0577] <= 174;
        weight_mem[16'h0578] <= 174;
        weight_mem[16'h0579] <= 181;
        weight_mem[16'h057A] <= 185;
        weight_mem[16'h057B] <= 184;
        weight_mem[16'h057C] <= 181;
        weight_mem[16'h057D] <= 179;
        weight_mem[16'h057E] <= 179;
        weight_mem[16'h057F] <= 179;
        weight_mem[16'h0580] <= 179;
        weight_mem[16'h0581] <= 179;
        weight_mem[16'h0582] <= 180;
        weight_mem[16'h0583] <= 180;
        weight_mem[16'h0584] <= 180;
        weight_mem[16'h0585] <= 181;
        weight_mem[16'h0586] <= 184;
        weight_mem[16'h0587] <= 186;
        weight_mem[16'h0588] <= 187;
        weight_mem[16'h0589] <= 195;
        weight_mem[16'h058A] <= 199;
        weight_mem[16'h058B] <= 186;
        weight_mem[16'h058C] <= 183;
        weight_mem[16'h058D] <= 191;
        weight_mem[16'h058E] <= 191;
        weight_mem[16'h058F] <= 185;
        weight_mem[16'h0590] <= 183;
        weight_mem[16'h0591] <= 183;
        weight_mem[16'h0592] <= 182;
        weight_mem[16'h0593] <= 182;
        weight_mem[16'h0594] <= 181;
        weight_mem[16'h0595] <= 179;
        weight_mem[16'h0596] <= 179;
        weight_mem[16'h0597] <= 179;
        weight_mem[16'h0598] <= 179;
        weight_mem[16'h0599] <= 179;
        weight_mem[16'h059A] <= 179;
        weight_mem[16'h059B] <= 179;
        weight_mem[16'h059C] <= 179;
        weight_mem[16'h059D] <= 180;
        weight_mem[16'h059E] <= 180;
        weight_mem[16'h059F] <= 181;
        weight_mem[16'h05A0] <= 180;
        weight_mem[16'h05A1] <= 180;
        weight_mem[16'h05A2] <= 181;
        weight_mem[16'h05A3] <= 178;
        weight_mem[16'h05A4] <= 178;
        weight_mem[16'h05A5] <= 179;
        weight_mem[16'h05A6] <= 180;
        weight_mem[16'h05A7] <= 179;
        weight_mem[16'h05A8] <= 180;
        weight_mem[16'h05A9] <= 180;
        weight_mem[16'h05AA] <= 180;
        weight_mem[16'h05AB] <= 179;
        weight_mem[16'h05AC] <= 179;
        weight_mem[16'h05AD] <= 179;
        weight_mem[16'h05AE] <= 179;
        weight_mem[16'h05AF] <= 179;

        // layer 1 neuron 3
        weight_mem[16'h0600] <= 252;
        weight_mem[16'h0601] <= 2;
        weight_mem[16'h0602] <= 9;
        weight_mem[16'h0603] <= 2;
        weight_mem[16'h0604] <= 250;
        weight_mem[16'h0605] <= 8;
        weight_mem[16'h0606] <= 10;
        weight_mem[16'h0607] <= 10;
        weight_mem[16'h0608] <= 252;
        weight_mem[16'h0609] <= 6;
        weight_mem[16'h060A] <= 248;
        weight_mem[16'h060B] <= 251;
        weight_mem[16'h060C] <= 11;
        weight_mem[16'h060D] <= 255;
        weight_mem[16'h060E] <= 249;
        weight_mem[16'h060F] <= 251;
        weight_mem[16'h0610] <= 244;
        weight_mem[16'h0611] <= 3;
        weight_mem[16'h0612] <= 246;
        weight_mem[16'h0613] <= 3;
        weight_mem[16'h0614] <= 255;
        weight_mem[16'h0615] <= 246;
        weight_mem[16'h0616] <= 254;
        weight_mem[16'h0617] <= 5;
        weight_mem[16'h0618] <= 250;
        weight_mem[16'h0619] <= 245;
        weight_mem[16'h061A] <= 1;
        weight_mem[16'h061B] <= 3;
        weight_mem[16'h061C] <= 6;
        weight_mem[16'h061D] <= 12;
        weight_mem[16'h061E] <= 247;
        weight_mem[16'h061F] <= 254;
        weight_mem[16'h0620] <= 12;
        weight_mem[16'h0621] <= 3;
        weight_mem[16'h0622] <= 13;
        weight_mem[16'h0623] <= 254;
        weight_mem[16'h0624] <= 9;
        weight_mem[16'h0625] <= 17;
        weight_mem[16'h0626] <= 5;
        weight_mem[16'h0627] <= 3;
        weight_mem[16'h0628] <= 5;
        weight_mem[16'h0629] <= 13;
        weight_mem[16'h062A] <= 9;
        weight_mem[16'h062B] <= 4;
        weight_mem[16'h062C] <= 11;
        weight_mem[16'h062D] <= 249;
        weight_mem[16'h062E] <= 248;
        weight_mem[16'h062F] <= 252;
        weight_mem[16'h0630] <= 246;
        weight_mem[16'h0631] <= 6;
        weight_mem[16'h0632] <= 2;
        weight_mem[16'h0633] <= 0;
        weight_mem[16'h0634] <= 253;
        weight_mem[16'h0635] <= 6;
        weight_mem[16'h0636] <= 12;
        weight_mem[16'h0637] <= 10;
        weight_mem[16'h0638] <= 13;
        weight_mem[16'h0639] <= 251;
        weight_mem[16'h063A] <= 11;
        weight_mem[16'h063B] <= 19;
        weight_mem[16'h063C] <= 8;
        weight_mem[16'h063D] <= 19;
        weight_mem[16'h063E] <= 22;
        weight_mem[16'h063F] <= 11;
        weight_mem[16'h0640] <= 23;
        weight_mem[16'h0641] <= 11;
        weight_mem[16'h0642] <= 9;
        weight_mem[16'h0643] <= 252;
        weight_mem[16'h0644] <= 253;
        weight_mem[16'h0645] <= 8;
        weight_mem[16'h0646] <= 245;
        weight_mem[16'h0647] <= 12;
        weight_mem[16'h0648] <= 253;
        weight_mem[16'h0649] <= 246;
        weight_mem[16'h064A] <= 3;
        weight_mem[16'h064B] <= 7;
        weight_mem[16'h064C] <= 2;
        weight_mem[16'h064D] <= 18;
        weight_mem[16'h064E] <= 7;
        weight_mem[16'h064F] <= 12;
        weight_mem[16'h0650] <= 10;
        weight_mem[16'h0651] <= 5;
        weight_mem[16'h0652] <= 255;
        weight_mem[16'h0653] <= 252;
        weight_mem[16'h0654] <= 23;
        weight_mem[16'h0655] <= 33;
        weight_mem[16'h0656] <= 42;
        weight_mem[16'h0657] <= 40;
        weight_mem[16'h0658] <= 30;
        weight_mem[16'h0659] <= 34;
        weight_mem[16'h065A] <= 33;
        weight_mem[16'h065B] <= 28;
        weight_mem[16'h065C] <= 22;
        weight_mem[16'h065D] <= 6;
        weight_mem[16'h065E] <= 252;
        weight_mem[16'h065F] <= 3;
        weight_mem[16'h0660] <= 245;
        weight_mem[16'h0661] <= 8;
        weight_mem[16'h0662] <= 254;
        weight_mem[16'h0663] <= 246;
        weight_mem[16'h0664] <= 14;
        weight_mem[16'h0665] <= 19;
        weight_mem[16'h0666] <= 22;
        weight_mem[16'h0667] <= 6;
        weight_mem[16'h0668] <= 252;
        weight_mem[16'h0669] <= 221;
        weight_mem[16'h066A] <= 202;
        weight_mem[16'h066B] <= 159;
        weight_mem[16'h066C] <= 133;
        weight_mem[16'h066D] <= 130;
        weight_mem[16'h066E] <= 155;
        weight_mem[16'h066F] <= 184;
        weight_mem[16'h0670] <= 222;
        weight_mem[16'h0671] <= 249;
        weight_mem[16'h0672] <= 31;
        weight_mem[16'h0673] <= 42;
        weight_mem[16'h0674] <= 31;
        weight_mem[16'h0675] <= 32;
        weight_mem[16'h0676] <= 16;
        weight_mem[16'h0677] <= 254;
        weight_mem[16'h0678] <= 2;
        weight_mem[16'h0679] <= 2;
        weight_mem[16'h067A] <= 4;
        weight_mem[16'h067B] <= 1;
        weight_mem[16'h067C] <= 254;
        weight_mem[16'h067D] <= 6;
        weight_mem[16'h067E] <= 10;
        weight_mem[16'h067F] <= 242;
        weight_mem[16'h0680] <= 216;
        weight_mem[16'h0681] <= 202;
        weight_mem[16'h0682] <= 185;
        weight_mem[16'h0683] <= 172;
        weight_mem[16'h0684] <= 128;
        weight_mem[16'h0685] <= 137;
        weight_mem[16'h0686] <= 172;
        weight_mem[16'h0687] <= 210;
        weight_mem[16'h0688] <= 237;
        weight_mem[16'h0689] <= 10;
        weight_mem[16'h068A] <= 4;
        weight_mem[16'h068B] <= 40;
        weight_mem[16'h068C] <= 28;
        weight_mem[16'h068D] <= 37;
        weight_mem[16'h068E] <= 3;
        weight_mem[16'h068F] <= 254;
        weight_mem[16'h0690] <= 4;
        weight_mem[16'h0691] <= 6;
        weight_mem[16'h0692] <= 249;
        weight_mem[16'h0693] <= 251;
        weight_mem[16'h0694] <= 3;
        weight_mem[16'h0695] <= 248;
        weight_mem[16'h0696] <= 252;
        weight_mem[16'h0697] <= 236;
        weight_mem[16'h0698] <= 217;
        weight_mem[16'h0699] <= 224;
        weight_mem[16'h069A] <= 234;
        weight_mem[16'h069B] <= 235;
        weight_mem[16'h069C] <= 228;
        weight_mem[16'h069D] <= 245;
        weight_mem[16'h069E] <= 241;
        weight_mem[16'h069F] <= 234;
        weight_mem[16'h06A0] <= 241;
        weight_mem[16'h06A1] <= 226;
        weight_mem[16'h06A2] <= 231;
        weight_mem[16'h06A3] <= 238;
        weight_mem[16'h06A4] <= 17;
        weight_mem[16'h06A5] <= 18;
        weight_mem[16'h06A6] <= 19;
        weight_mem[16'h06A7] <= 5;
        weight_mem[16'h06A8] <= 9;
        weight_mem[16'h06A9] <= 7;
        weight_mem[16'h06AA] <= 254;
        weight_mem[16'h06AB] <= 247;
        weight_mem[16'h06AC] <= 237;
        weight_mem[16'h06AD] <= 225;
        weight_mem[16'h06AE] <= 220;
        weight_mem[16'h06AF] <= 238;
        weight_mem[16'h06B0] <= 244;
        weight_mem[16'h06B1] <= 243;
        weight_mem[16'h06B2] <= 28;
        weight_mem[16'h06B3] <= 43;
        weight_mem[16'h06B4] <= 56;
        weight_mem[16'h06B5] <= 43;
        weight_mem[16'h06B6] <= 251;
        weight_mem[16'h06B7] <= 193;
        weight_mem[16'h06B8] <= 192;
        weight_mem[16'h06B9] <= 196;
        weight_mem[16'h06BA] <= 202;
        weight_mem[16'h06BB] <= 211;
        weight_mem[16'h06BC] <= 253;
        weight_mem[16'h06BD] <= 2;
        weight_mem[16'h06BE] <= 254;
        weight_mem[16'h06BF] <= 12;
        weight_mem[16'h06C0] <= 254;
        weight_mem[16'h06C1] <= 11;
        weight_mem[16'h06C2] <= 5;
        weight_mem[16'h06C3] <= 251;
        weight_mem[16'h06C4] <= 236;
        weight_mem[16'h06C5] <= 221;
        weight_mem[16'h06C6] <= 216;
        weight_mem[16'h06C7] <= 0;
        weight_mem[16'h06C8] <= 8;
        weight_mem[16'h06C9] <= 45;
        weight_mem[16'h06CA] <= 93;
        weight_mem[16'h06CB] <= 84;
        weight_mem[16'h06CC] <= 38;
        weight_mem[16'h06CD] <= 12;
        weight_mem[16'h06CE] <= 218;
        weight_mem[16'h06CF] <= 205;
        weight_mem[16'h06D0] <= 215;
        weight_mem[16'h06D1] <= 222;
        weight_mem[16'h06D2] <= 216;
        weight_mem[16'h06D3] <= 213;
        weight_mem[16'h06D4] <= 246;
        weight_mem[16'h06D5] <= 10;
        weight_mem[16'h06D6] <= 3;
        weight_mem[16'h06D7] <= 6;
        weight_mem[16'h06D8] <= 1;
        weight_mem[16'h06D9] <= 244;
        weight_mem[16'h06DA] <= 249;
        weight_mem[16'h06DB] <= 243;
        weight_mem[16'h06DC] <= 245;
        weight_mem[16'h06DD] <= 227;
        weight_mem[16'h06DE] <= 245;
        weight_mem[16'h06DF] <= 9;
        weight_mem[16'h06E0] <= 6;
        weight_mem[16'h06E1] <= 17;
        weight_mem[16'h06E2] <= 40;
        weight_mem[16'h06E3] <= 41;
        weight_mem[16'h06E4] <= 47;
        weight_mem[16'h06E5] <= 13;
        weight_mem[16'h06E6] <= 225;
        weight_mem[16'h06E7] <= 245;
        weight_mem[16'h06E8] <= 249;
        weight_mem[16'h06E9] <= 238;
        weight_mem[16'h06EA] <= 244;
        weight_mem[16'h06EB] <= 3;
        weight_mem[16'h06EC] <= 5;
        weight_mem[16'h06ED] <= 12;
        weight_mem[16'h06EE] <= 248;
        weight_mem[16'h06EF] <= 255;
        weight_mem[16'h06F0] <= 0;
        weight_mem[16'h06F1] <= 253;
        weight_mem[16'h06F2] <= 0;
        weight_mem[16'h06F3] <= 6;
        weight_mem[16'h06F4] <= 4;
        weight_mem[16'h06F5] <= 12;
        weight_mem[16'h06F6] <= 250;
        weight_mem[16'h06F7] <= 246;
        weight_mem[16'h06F8] <= 226;
        weight_mem[16'h06F9] <= 211;
        weight_mem[16'h06FA] <= 250;
        weight_mem[16'h06FB] <= 74;
        weight_mem[16'h06FC] <= 115;
        weight_mem[16'h06FD] <= 57;
        weight_mem[16'h06FE] <= 4;
        weight_mem[16'h06FF] <= 249;
        weight_mem[16'h0700] <= 11;
        weight_mem[16'h0701] <= 4;
        weight_mem[16'h0702] <= 12;
        weight_mem[16'h0703] <= 11;
        weight_mem[16'h0704] <= 22;
        weight_mem[16'h0705] <= 1;
        weight_mem[16'h0706] <= 254;
        weight_mem[16'h0707] <= 4;
        weight_mem[16'h0708] <= 248;
        weight_mem[16'h0709] <= 5;
        weight_mem[16'h070A] <= 249;
        weight_mem[16'h070B] <= 3;
        weight_mem[16'h070C] <= 17;
        weight_mem[16'h070D] <= 20;
        weight_mem[16'h070E] <= 17;
        weight_mem[16'h070F] <= 241;
        weight_mem[16'h0710] <= 221;
        weight_mem[16'h0711] <= 215;
        weight_mem[16'h0712] <= 242;
        weight_mem[16'h0713] <= 58;
        weight_mem[16'h0714] <= 72;
        weight_mem[16'h0715] <= 35;
        weight_mem[16'h0716] <= 13;
        weight_mem[16'h0717] <= 247;
        weight_mem[16'h0718] <= 5;
        weight_mem[16'h0719] <= 8;
        weight_mem[16'h071A] <= 19;
        weight_mem[16'h071B] <= 32;
        weight_mem[16'h071C] <= 31;
        weight_mem[16'h071D] <= 18;
        weight_mem[16'h071E] <= 249;
        weight_mem[16'h071F] <= 250;
        weight_mem[16'h0720] <= 3;
        weight_mem[16'h0721] <= 250;
        weight_mem[16'h0722] <= 254;
        weight_mem[16'h0723] <= 11;
        weight_mem[16'h0724] <= 24;
        weight_mem[16'h0725] <= 39;
        weight_mem[16'h0726] <= 38;
        weight_mem[16'h0727] <= 15;
        weight_mem[16'h0728] <= 21;
        weight_mem[16'h0729] <= 254;
        weight_mem[16'h072A] <= 34;
        weight_mem[16'h072B] <= 30;
        weight_mem[16'h072C] <= 39;
        weight_mem[16'h072D] <= 37;
        weight_mem[16'h072E] <= 19;
        weight_mem[16'h072F] <= 11;
        weight_mem[16'h0730] <= 250;
        weight_mem[16'h0731] <= 255;
        weight_mem[16'h0732] <= 30;
        weight_mem[16'h0733] <= 32;
        weight_mem[16'h0734] <= 11;
        weight_mem[16'h0735] <= 12;
        weight_mem[16'h0736] <= 8;
        weight_mem[16'h0737] <= 249;
        weight_mem[16'h0738] <= 245;
        weight_mem[16'h0739] <= 10;
        weight_mem[16'h073A] <= 248;
        weight_mem[16'h073B] <= 14;
        weight_mem[16'h073C] <= 11;
        weight_mem[16'h073D] <= 21;
        weight_mem[16'h073E] <= 54;
        weight_mem[16'h073F] <= 39;
        weight_mem[16'h0740] <= 43;
        weight_mem[16'h0741] <= 29;
        weight_mem[16'h0742] <= 38;
        weight_mem[16'h0743] <= 29;
        weight_mem[16'h0744] <= 32;
        weight_mem[16'h0745] <= 20;
        weight_mem[16'h0746] <= 25;
        weight_mem[16'h0747] <= 33;
        weight_mem[16'h0748] <= 28;
        weight_mem[16'h0749] <= 33;
        weight_mem[16'h074A] <= 31;
        weight_mem[16'h074B] <= 24;
        weight_mem[16'h074C] <= 19;
        weight_mem[16'h074D] <= 5;
        weight_mem[16'h074E] <= 254;
        weight_mem[16'h074F] <= 252;
        weight_mem[16'h0750] <= 255;
        weight_mem[16'h0751] <= 254;
        weight_mem[16'h0752] <= 253;
        weight_mem[16'h0753] <= 13;
        weight_mem[16'h0754] <= 1;
        weight_mem[16'h0755] <= 7;
        weight_mem[16'h0756] <= 7;
        weight_mem[16'h0757] <= 16;
        weight_mem[16'h0758] <= 4;
        weight_mem[16'h0759] <= 18;
        weight_mem[16'h075A] <= 1;
        weight_mem[16'h075B] <= 17;
        weight_mem[16'h075C] <= 6;
        weight_mem[16'h075D] <= 31;
        weight_mem[16'h075E] <= 37;
        weight_mem[16'h075F] <= 41;
        weight_mem[16'h0760] <= 57;
        weight_mem[16'h0761] <= 27;
        weight_mem[16'h0762] <= 20;
        weight_mem[16'h0763] <= 0;
        weight_mem[16'h0764] <= 4;
        weight_mem[16'h0765] <= 248;
        weight_mem[16'h0766] <= 9;
        weight_mem[16'h0767] <= 7;
        weight_mem[16'h0768] <= 254;
        weight_mem[16'h0769] <= 252;
        weight_mem[16'h076A] <= 253;
        weight_mem[16'h076B] <= 8;
        weight_mem[16'h076C] <= 244;
        weight_mem[16'h076D] <= 246;
        weight_mem[16'h076E] <= 243;
        weight_mem[16'h076F] <= 239;
        weight_mem[16'h0770] <= 235;
        weight_mem[16'h0771] <= 2;
        weight_mem[16'h0772] <= 7;
        weight_mem[16'h0773] <= 10;
        weight_mem[16'h0774] <= 43;
        weight_mem[16'h0775] <= 31;
        weight_mem[16'h0776] <= 14;
        weight_mem[16'h0777] <= 0;
        weight_mem[16'h0778] <= 255;
        weight_mem[16'h0779] <= 245;
        weight_mem[16'h077A] <= 0;
        weight_mem[16'h077B] <= 254;
        weight_mem[16'h077C] <= 255;
        weight_mem[16'h077D] <= 5;
        weight_mem[16'h077E] <= 254;
        weight_mem[16'h077F] <= 7;
        weight_mem[16'h0780] <= 3;
        weight_mem[16'h0781] <= 12;
        weight_mem[16'h0782] <= 8;
        weight_mem[16'h0783] <= 1;
        weight_mem[16'h0784] <= 1;
        weight_mem[16'h0785] <= 245;
        weight_mem[16'h0786] <= 231;
        weight_mem[16'h0787] <= 218;
        weight_mem[16'h0788] <= 225;
        weight_mem[16'h0789] <= 213;
        weight_mem[16'h078A] <= 222;
        weight_mem[16'h078B] <= 229;
        weight_mem[16'h078C] <= 219;
        weight_mem[16'h078D] <= 236;
        weight_mem[16'h078E] <= 220;
        weight_mem[16'h078F] <= 215;
        weight_mem[16'h0790] <= 236;
        weight_mem[16'h0791] <= 239;
        weight_mem[16'h0792] <= 247;
        weight_mem[16'h0793] <= 251;
        weight_mem[16'h0794] <= 253;
        weight_mem[16'h0795] <= 252;
        weight_mem[16'h0796] <= 249;
        weight_mem[16'h0797] <= 2;
        weight_mem[16'h0798] <= 252;
        weight_mem[16'h0799] <= 1;
        weight_mem[16'h079A] <= 3;
        weight_mem[16'h079B] <= 5;
        weight_mem[16'h079C] <= 248;
        weight_mem[16'h079D] <= 255;
        weight_mem[16'h079E] <= 240;
        weight_mem[16'h079F] <= 247;
        weight_mem[16'h07A0] <= 252;
        weight_mem[16'h07A1] <= 250;
        weight_mem[16'h07A2] <= 244;
        weight_mem[16'h07A3] <= 233;
        weight_mem[16'h07A4] <= 228;
        weight_mem[16'h07A5] <= 241;
        weight_mem[16'h07A6] <= 248;
        weight_mem[16'h07A7] <= 243;
        weight_mem[16'h07A8] <= 246;
        weight_mem[16'h07A9] <= 242;
        weight_mem[16'h07AA] <= 248;
        weight_mem[16'h07AB] <= 1;
        weight_mem[16'h07AC] <= 253;
        weight_mem[16'h07AD] <= 5;
        weight_mem[16'h07AE] <= 8;
        weight_mem[16'h07AF] <= 11;

        // layer 1 neuron 4
        weight_mem[16'h0800] <= 253;
        weight_mem[16'h0801] <= 248;
        weight_mem[16'h0802] <= 7;
        weight_mem[16'h0803] <= 0;
        weight_mem[16'h0804] <= 6;
        weight_mem[16'h0805] <= 254;
        weight_mem[16'h0806] <= 251;
        weight_mem[16'h0807] <= 8;
        weight_mem[16'h0808] <= 255;
        weight_mem[16'h0809] <= 8;
        weight_mem[16'h080A] <= 3;
        weight_mem[16'h080B] <= 8;
        weight_mem[16'h080C] <= 8;
        weight_mem[16'h080D] <= 3;
        weight_mem[16'h080E] <= 7;
        weight_mem[16'h080F] <= 250;
        weight_mem[16'h0810] <= 0;
        weight_mem[16'h0811] <= 10;
        weight_mem[16'h0812] <= 3;
        weight_mem[16'h0813] <= 1;
        weight_mem[16'h0814] <= 255;
        weight_mem[16'h0815] <= 249;
        weight_mem[16'h0816] <= 254;
        weight_mem[16'h0817] <= 1;
        weight_mem[16'h0818] <= 6;
        weight_mem[16'h0819] <= 3;
        weight_mem[16'h081A] <= 4;
        weight_mem[16'h081B] <= 252;
        weight_mem[16'h081C] <= 255;
        weight_mem[16'h081D] <= 252;
        weight_mem[16'h081E] <= 9;
        weight_mem[16'h081F] <= 1;
        weight_mem[16'h0820] <= 248;
        weight_mem[16'h0821] <= 3;
        weight_mem[16'h0822] <= 0;
        weight_mem[16'h0823] <= 5;
        weight_mem[16'h0824] <= 251;
        weight_mem[16'h0825] <= 11;
        weight_mem[16'h0826] <= 9;
        weight_mem[16'h0827] <= 5;
        weight_mem[16'h0828] <= 1;
        weight_mem[16'h0829] <= 9;
        weight_mem[16'h082A] <= 251;
        weight_mem[16'h082B] <= 7;
        weight_mem[16'h082C] <= 3;
        weight_mem[16'h082D] <= 10;
        weight_mem[16'h082E] <= 253;
        weight_mem[16'h082F] <= 254;
        weight_mem[16'h0830] <= 1;
        weight_mem[16'h0831] <= 8;
        weight_mem[16'h0832] <= 5;
        weight_mem[16'h0833] <= 250;
        weight_mem[16'h0834] <= 248;
        weight_mem[16'h0835] <= 255;
        weight_mem[16'h0836] <= 252;
        weight_mem[16'h0837] <= 238;
        weight_mem[16'h0838] <= 239;
        weight_mem[16'h0839] <= 219;
        weight_mem[16'h083A] <= 217;
        weight_mem[16'h083B] <= 222;
        weight_mem[16'h083C] <= 224;
        weight_mem[16'h083D] <= 235;
        weight_mem[16'h083E] <= 242;
        weight_mem[16'h083F] <= 0;
        weight_mem[16'h0840] <= 7;
        weight_mem[16'h0841] <= 18;
        weight_mem[16'h0842] <= 12;
        weight_mem[16'h0843] <= 1;
        weight_mem[16'h0844] <= 255;
        weight_mem[16'h0845] <= 10;
        weight_mem[16'h0846] <= 3;
        weight_mem[16'h0847] <= 254;
        weight_mem[16'h0848] <= 253;
        weight_mem[16'h0849] <= 254;
        weight_mem[16'h084A] <= 252;
        weight_mem[16'h084B] <= 244;
        weight_mem[16'h084C] <= 250;
        weight_mem[16'h084D] <= 232;
        weight_mem[16'h084E] <= 244;
        weight_mem[16'h084F] <= 228;
        weight_mem[16'h0850] <= 232;
        weight_mem[16'h0851] <= 220;
        weight_mem[16'h0852] <= 219;
        weight_mem[16'h0853] <= 245;
        weight_mem[16'h0854] <= 246;
        weight_mem[16'h0855] <= 2;
        weight_mem[16'h0856] <= 244;
        weight_mem[16'h0857] <= 251;
        weight_mem[16'h0858] <= 6;
        weight_mem[16'h0859] <= 7;
        weight_mem[16'h085A] <= 5;
        weight_mem[16'h085B] <= 13;
        weight_mem[16'h085C] <= 252;
        weight_mem[16'h085D] <= 253;
        weight_mem[16'h085E] <= 253;
        weight_mem[16'h085F] <= 7;
        weight_mem[16'h0860] <= 249;
        weight_mem[16'h0861] <= 251;
        weight_mem[16'h0862] <= 250;
        weight_mem[16'h0863] <= 243;
        weight_mem[16'h0864] <= 239;
        weight_mem[16'h0865] <= 239;
        weight_mem[16'h0866] <= 246;
        weight_mem[16'h0867] <= 0;
        weight_mem[16'h0868] <= 248;
        weight_mem[16'h0869] <= 250;
        weight_mem[16'h086A] <= 250;
        weight_mem[16'h086B] <= 231;
        weight_mem[16'h086C] <= 230;
        weight_mem[16'h086D] <= 247;
        weight_mem[16'h086E] <= 238;
        weight_mem[16'h086F] <= 236;
        weight_mem[16'h0870] <= 248;
        weight_mem[16'h0871] <= 244;
        weight_mem[16'h0872] <= 251;
        weight_mem[16'h0873] <= 254;
        weight_mem[16'h0874] <= 5;
        weight_mem[16'h0875] <= 1;
        weight_mem[16'h0876] <= 248;
        weight_mem[16'h0877] <= 253;
        weight_mem[16'h0878] <= 5;
        weight_mem[16'h0879] <= 250;
        weight_mem[16'h087A] <= 252;
        weight_mem[16'h087B] <= 244;
        weight_mem[16'h087C] <= 242;
        weight_mem[16'h087D] <= 244;
        weight_mem[16'h087E] <= 13;
        weight_mem[16'h087F] <= 8;
        weight_mem[16'h0880] <= 17;
        weight_mem[16'h0881] <= 1;
        weight_mem[16'h0882] <= 246;
        weight_mem[16'h0883] <= 223;
        weight_mem[16'h0884] <= 216;
        weight_mem[16'h0885] <= 218;
        weight_mem[16'h0886] <= 246;
        weight_mem[16'h0887] <= 8;
        weight_mem[16'h0888] <= 8;
        weight_mem[16'h0889] <= 253;
        weight_mem[16'h088A] <= 253;
        weight_mem[16'h088B] <= 8;
        weight_mem[16'h088C] <= 9;
        weight_mem[16'h088D] <= 251;
        weight_mem[16'h088E] <= 2;
        weight_mem[16'h088F] <= 248;
        weight_mem[16'h0890] <= 1;
        weight_mem[16'h0891] <= 253;
        weight_mem[16'h0892] <= 252;
        weight_mem[16'h0893] <= 252;
        weight_mem[16'h0894] <= 4;
        weight_mem[16'h0895] <= 4;
        weight_mem[16'h0896] <= 19;
        weight_mem[16'h0897] <= 29;
        weight_mem[16'h0898] <= 30;
        weight_mem[16'h0899] <= 27;
        weight_mem[16'h089A] <= 36;
        weight_mem[16'h089B] <= 19;
        weight_mem[16'h089C] <= 251;
        weight_mem[16'h089D] <= 255;
        weight_mem[16'h089E] <= 18;
        weight_mem[16'h089F] <= 15;
        weight_mem[16'h08A0] <= 20;
        weight_mem[16'h08A1] <= 10;
        weight_mem[16'h08A2] <= 18;
        weight_mem[16'h08A3] <= 16;
        weight_mem[16'h08A4] <= 14;
        weight_mem[16'h08A5] <= 255;
        weight_mem[16'h08A6] <= 9;
        weight_mem[16'h08A7] <= 8;
        weight_mem[16'h08A8] <= 0;
        weight_mem[16'h08A9] <= 0;
        weight_mem[16'h08AA] <= 0;
        weight_mem[16'h08AB] <= 9;
        weight_mem[16'h08AC] <= 14;
        weight_mem[16'h08AD] <= 35;
        weight_mem[16'h08AE] <= 46;
        weight_mem[16'h08AF] <= 35;
        weight_mem[16'h08B0] <= 23;
        weight_mem[16'h08B1] <= 13;
        weight_mem[16'h08B2] <= 249;
        weight_mem[16'h08B3] <= 225;
        weight_mem[16'h08B4] <= 231;
        weight_mem[16'h08B5] <= 0;
        weight_mem[16'h08B6] <= 12;
        weight_mem[16'h08B7] <= 243;
        weight_mem[16'h08B8] <= 1;
        weight_mem[16'h08B9] <= 15;
        weight_mem[16'h08BA] <= 43;
        weight_mem[16'h08BB] <= 20;
        weight_mem[16'h08BC] <= 8;
        weight_mem[16'h08BD] <= 253;
        weight_mem[16'h08BE] <= 10;
        weight_mem[16'h08BF] <= 251;
        weight_mem[16'h08C0] <= 1;
        weight_mem[16'h08C1] <= 250;
        weight_mem[16'h08C2] <= 254;
        weight_mem[16'h08C3] <= 1;
        weight_mem[16'h08C4] <= 14;
        weight_mem[16'h08C5] <= 27;
        weight_mem[16'h08C6] <= 23;
        weight_mem[16'h08C7] <= 12;
        weight_mem[16'h08C8] <= 241;
        weight_mem[16'h08C9] <= 241;
        weight_mem[16'h08CA] <= 232;
        weight_mem[16'h08CB] <= 221;
        weight_mem[16'h08CC] <= 227;
        weight_mem[16'h08CD] <= 13;
        weight_mem[16'h08CE] <= 254;
        weight_mem[16'h08CF] <= 242;
        weight_mem[16'h08D0] <= 7;
        weight_mem[16'h08D1] <= 26;
        weight_mem[16'h08D2] <= 44;
        weight_mem[16'h08D3] <= 27;
        weight_mem[16'h08D4] <= 24;
        weight_mem[16'h08D5] <= 7;
        weight_mem[16'h08D6] <= 9;
        weight_mem[16'h08D7] <= 250;
        weight_mem[16'h08D8] <= 0;
        weight_mem[16'h08D9] <= 0;
        weight_mem[16'h08DA] <= 251;
        weight_mem[16'h08DB] <= 3;
        weight_mem[16'h08DC] <= 11;
        weight_mem[16'h08DD] <= 23;
        weight_mem[16'h08DE] <= 28;
        weight_mem[16'h08DF] <= 18;
        weight_mem[16'h08E0] <= 244;
        weight_mem[16'h08E1] <= 244;
        weight_mem[16'h08E2] <= 247;
        weight_mem[16'h08E3] <= 225;
        weight_mem[16'h08E4] <= 239;
        weight_mem[16'h08E5] <= 4;
        weight_mem[16'h08E6] <= 250;
        weight_mem[16'h08E7] <= 252;
        weight_mem[16'h08E8] <= 255;
        weight_mem[16'h08E9] <= 254;
        weight_mem[16'h08EA] <= 1;
        weight_mem[16'h08EB] <= 7;
        weight_mem[16'h08EC] <= 14;
        weight_mem[16'h08ED] <= 3;
        weight_mem[16'h08EE] <= 8;
        weight_mem[16'h08EF] <= 253;
        weight_mem[16'h08F0] <= 2;
        weight_mem[16'h08F1] <= 7;
        weight_mem[16'h08F2] <= 2;
        weight_mem[16'h08F3] <= 252;
        weight_mem[16'h08F4] <= 9;
        weight_mem[16'h08F5] <= 38;
        weight_mem[16'h08F6] <= 56;
        weight_mem[16'h08F7] <= 81;
        weight_mem[16'h08F8] <= 69;
        weight_mem[16'h08F9] <= 45;
        weight_mem[16'h08FA] <= 16;
        weight_mem[16'h08FB] <= 6;
        weight_mem[16'h08FC] <= 33;
        weight_mem[16'h08FD] <= 15;
        weight_mem[16'h08FE] <= 5;
        weight_mem[16'h08FF] <= 4;
        weight_mem[16'h0900] <= 240;
        weight_mem[16'h0901] <= 222;
        weight_mem[16'h0902] <= 231;
        weight_mem[16'h0903] <= 232;
        weight_mem[16'h0904] <= 255;
        weight_mem[16'h0905] <= 9;
        weight_mem[16'h0906] <= 2;
        weight_mem[16'h0907] <= 248;
        weight_mem[16'h0908] <= 8;
        weight_mem[16'h0909] <= 8;
        weight_mem[16'h090A] <= 249;
        weight_mem[16'h090B] <= 244;
        weight_mem[16'h090C] <= 234;
        weight_mem[16'h090D] <= 19;
        weight_mem[16'h090E] <= 56;
        weight_mem[16'h090F] <= 100;
        weight_mem[16'h0910] <= 127;
        weight_mem[16'h0911] <= 124;
        weight_mem[16'h0912] <= 124;
        weight_mem[16'h0913] <= 86;
        weight_mem[16'h0914] <= 43;
        weight_mem[16'h0915] <= 253;
        weight_mem[16'h0916] <= 243;
        weight_mem[16'h0917] <= 247;
        weight_mem[16'h0918] <= 225;
        weight_mem[16'h0919] <= 230;
        weight_mem[16'h091A] <= 206;
        weight_mem[16'h091B] <= 224;
        weight_mem[16'h091C] <= 250;
        weight_mem[16'h091D] <= 3;
        weight_mem[16'h091E] <= 0;
        weight_mem[16'h091F] <= 251;
        weight_mem[16'h0920] <= 253;
        weight_mem[16'h0921] <= 255;
        weight_mem[16'h0922] <= 253;
        weight_mem[16'h0923] <= 227;
        weight_mem[16'h0924] <= 221;
        weight_mem[16'h0925] <= 236;
        weight_mem[16'h0926] <= 5;
        weight_mem[16'h0927] <= 17;
        weight_mem[16'h0928] <= 37;
        weight_mem[16'h0929] <= 47;
        weight_mem[16'h092A] <= 66;
        weight_mem[16'h092B] <= 39;
        weight_mem[16'h092C] <= 250;
        weight_mem[16'h092D] <= 233;
        weight_mem[16'h092E] <= 229;
        weight_mem[16'h092F] <= 234;
        weight_mem[16'h0930] <= 228;
        weight_mem[16'h0931] <= 216;
        weight_mem[16'h0932] <= 222;
        weight_mem[16'h0933] <= 232;
        weight_mem[16'h0934] <= 5;
        weight_mem[16'h0935] <= 7;
        weight_mem[16'h0936] <= 6;
        weight_mem[16'h0937] <= 254;
        weight_mem[16'h0938] <= 9;
        weight_mem[16'h0939] <= 255;
        weight_mem[16'h093A] <= 244;
        weight_mem[16'h093B] <= 238;
        weight_mem[16'h093C] <= 233;
        weight_mem[16'h093D] <= 224;
        weight_mem[16'h093E] <= 232;
        weight_mem[16'h093F] <= 228;
        weight_mem[16'h0940] <= 235;
        weight_mem[16'h0941] <= 242;
        weight_mem[16'h0942] <= 235;
        weight_mem[16'h0943] <= 233;
        weight_mem[16'h0944] <= 232;
        weight_mem[16'h0945] <= 238;
        weight_mem[16'h0946] <= 249;
        weight_mem[16'h0947] <= 243;
        weight_mem[16'h0948] <= 236;
        weight_mem[16'h0949] <= 241;
        weight_mem[16'h094A] <= 254;
        weight_mem[16'h094B] <= 253;
        weight_mem[16'h094C] <= 15;
        weight_mem[16'h094D] <= 5;
        weight_mem[16'h094E] <= 249;
        weight_mem[16'h094F] <= 254;
        weight_mem[16'h0950] <= 4;
        weight_mem[16'h0951] <= 4;
        weight_mem[16'h0952] <= 2;
        weight_mem[16'h0953] <= 243;
        weight_mem[16'h0954] <= 244;
        weight_mem[16'h0955] <= 239;
        weight_mem[16'h0956] <= 245;
        weight_mem[16'h0957] <= 244;
        weight_mem[16'h0958] <= 244;
        weight_mem[16'h0959] <= 231;
        weight_mem[16'h095A] <= 248;
        weight_mem[16'h095B] <= 250;
        weight_mem[16'h095C] <= 13;
        weight_mem[16'h095D] <= 14;
        weight_mem[16'h095E] <= 6;
        weight_mem[16'h095F] <= 0;
        weight_mem[16'h0960] <= 8;
        weight_mem[16'h0961] <= 254;
        weight_mem[16'h0962] <= 15;
        weight_mem[16'h0963] <= 6;
        weight_mem[16'h0964] <= 251;
        weight_mem[16'h0965] <= 9;
        weight_mem[16'h0966] <= 1;
        weight_mem[16'h0967] <= 2;
        weight_mem[16'h0968] <= 2;
        weight_mem[16'h0969] <= 250;
        weight_mem[16'h096A] <= 252;
        weight_mem[16'h096B] <= 241;
        weight_mem[16'h096C] <= 233;
        weight_mem[16'h096D] <= 233;
        weight_mem[16'h096E] <= 218;
        weight_mem[16'h096F] <= 233;
        weight_mem[16'h0970] <= 235;
        weight_mem[16'h0971] <= 231;
        weight_mem[16'h0972] <= 245;
        weight_mem[16'h0973] <= 245;
        weight_mem[16'h0974] <= 0;
        weight_mem[16'h0975] <= 16;
        weight_mem[16'h0976] <= 5;
        weight_mem[16'h0977] <= 19;
        weight_mem[16'h0978] <= 16;
        weight_mem[16'h0979] <= 14;
        weight_mem[16'h097A] <= 4;
        weight_mem[16'h097B] <= 8;
        weight_mem[16'h097C] <= 5;
        weight_mem[16'h097D] <= 6;
        weight_mem[16'h097E] <= 7;
        weight_mem[16'h097F] <= 5;
        weight_mem[16'h0980] <= 6;
        weight_mem[16'h0981] <= 5;
        weight_mem[16'h0982] <= 250;
        weight_mem[16'h0983] <= 250;
        weight_mem[16'h0984] <= 244;
        weight_mem[16'h0985] <= 255;
        weight_mem[16'h0986] <= 249;
        weight_mem[16'h0987] <= 229;
        weight_mem[16'h0988] <= 228;
        weight_mem[16'h0989] <= 225;
        weight_mem[16'h098A] <= 234;
        weight_mem[16'h098B] <= 223;
        weight_mem[16'h098C] <= 243;
        weight_mem[16'h098D] <= 251;
        weight_mem[16'h098E] <= 246;
        weight_mem[16'h098F] <= 250;
        weight_mem[16'h0990] <= 248;
        weight_mem[16'h0991] <= 253;
        weight_mem[16'h0992] <= 254;
        weight_mem[16'h0993] <= 9;
        weight_mem[16'h0994] <= 0;
        weight_mem[16'h0995] <= 249;
        weight_mem[16'h0996] <= 1;
        weight_mem[16'h0997] <= 9;
        weight_mem[16'h0998] <= 6;
        weight_mem[16'h0999] <= 1;
        weight_mem[16'h099A] <= 251;
        weight_mem[16'h099B] <= 7;
        weight_mem[16'h099C] <= 9;
        weight_mem[16'h099D] <= 254;
        weight_mem[16'h099E] <= 253;
        weight_mem[16'h099F] <= 5;
        weight_mem[16'h09A0] <= 3;
        weight_mem[16'h09A1] <= 1;
        weight_mem[16'h09A2] <= 4;
        weight_mem[16'h09A3] <= 3;
        weight_mem[16'h09A4] <= 4;
        weight_mem[16'h09A5] <= 5;
        weight_mem[16'h09A6] <= 247;
        weight_mem[16'h09A7] <= 7;
        weight_mem[16'h09A8] <= 250;
        weight_mem[16'h09A9] <= 6;
        weight_mem[16'h09AA] <= 248;
        weight_mem[16'h09AB] <= 9;
        weight_mem[16'h09AC] <= 252;
        weight_mem[16'h09AD] <= 7;
        weight_mem[16'h09AE] <= 6;
        weight_mem[16'h09AF] <= 9;

        // layer 1 neuron 5
        weight_mem[16'h0A00] <= 0;
        weight_mem[16'h0A01] <= 0;
        weight_mem[16'h0A02] <= 0;
        weight_mem[16'h0A03] <= 0;
        weight_mem[16'h0A04] <= 0;
        weight_mem[16'h0A05] <= 0;
        weight_mem[16'h0A06] <= 0;
        weight_mem[16'h0A07] <= 0;
        weight_mem[16'h0A08] <= 0;
        weight_mem[16'h0A09] <= 0;
        weight_mem[16'h0A0A] <= 0;
        weight_mem[16'h0A0B] <= 0;
        weight_mem[16'h0A0C] <= 0;
        weight_mem[16'h0A0D] <= 0;
        weight_mem[16'h0A0E] <= 0;
        weight_mem[16'h0A0F] <= 0;
        weight_mem[16'h0A10] <= 0;
        weight_mem[16'h0A11] <= 0;
        weight_mem[16'h0A12] <= 0;
        weight_mem[16'h0A13] <= 0;
        weight_mem[16'h0A14] <= 0;
        weight_mem[16'h0A15] <= 0;
        weight_mem[16'h0A16] <= 0;
        weight_mem[16'h0A17] <= 0;
        weight_mem[16'h0A18] <= 0;
        weight_mem[16'h0A19] <= 0;
        weight_mem[16'h0A1A] <= 0;
        weight_mem[16'h0A1B] <= 0;
        weight_mem[16'h0A1C] <= 0;
        weight_mem[16'h0A1D] <= 0;
        weight_mem[16'h0A1E] <= 0;
        weight_mem[16'h0A1F] <= 0;
        weight_mem[16'h0A20] <= 0;
        weight_mem[16'h0A21] <= 0;
        weight_mem[16'h0A22] <= 0;
        weight_mem[16'h0A23] <= 0;
        weight_mem[16'h0A24] <= 0;
        weight_mem[16'h0A25] <= 0;
        weight_mem[16'h0A26] <= 0;
        weight_mem[16'h0A27] <= 0;
        weight_mem[16'h0A28] <= 0;
        weight_mem[16'h0A29] <= 0;
        weight_mem[16'h0A2A] <= 0;
        weight_mem[16'h0A2B] <= 0;
        weight_mem[16'h0A2C] <= 0;
        weight_mem[16'h0A2D] <= 0;
        weight_mem[16'h0A2E] <= 0;
        weight_mem[16'h0A2F] <= 0;
        weight_mem[16'h0A30] <= 0;
        weight_mem[16'h0A31] <= 0;
        weight_mem[16'h0A32] <= 0;
        weight_mem[16'h0A33] <= 0;
        weight_mem[16'h0A34] <= 0;
        weight_mem[16'h0A35] <= 0;
        weight_mem[16'h0A36] <= 0;
        weight_mem[16'h0A37] <= 0;
        weight_mem[16'h0A38] <= 0;
        weight_mem[16'h0A39] <= 0;
        weight_mem[16'h0A3A] <= 0;
        weight_mem[16'h0A3B] <= 0;
        weight_mem[16'h0A3C] <= 0;
        weight_mem[16'h0A3D] <= 0;
        weight_mem[16'h0A3E] <= 0;
        weight_mem[16'h0A3F] <= 0;
        weight_mem[16'h0A40] <= 0;
        weight_mem[16'h0A41] <= 0;
        weight_mem[16'h0A42] <= 0;
        weight_mem[16'h0A43] <= 0;
        weight_mem[16'h0A44] <= 0;
        weight_mem[16'h0A45] <= 0;
        weight_mem[16'h0A46] <= 0;
        weight_mem[16'h0A47] <= 0;
        weight_mem[16'h0A48] <= 0;
        weight_mem[16'h0A49] <= 0;
        weight_mem[16'h0A4A] <= 0;
        weight_mem[16'h0A4B] <= 0;
        weight_mem[16'h0A4C] <= 0;
        weight_mem[16'h0A4D] <= 0;
        weight_mem[16'h0A4E] <= 0;
        weight_mem[16'h0A4F] <= 0;
        weight_mem[16'h0A50] <= 0;
        weight_mem[16'h0A51] <= 0;
        weight_mem[16'h0A52] <= 1;
        weight_mem[16'h0A53] <= 0;
        weight_mem[16'h0A54] <= 0;
        weight_mem[16'h0A55] <= 0;
        weight_mem[16'h0A56] <= 0;
        weight_mem[16'h0A57] <= 0;
        weight_mem[16'h0A58] <= 0;
        weight_mem[16'h0A59] <= 0;
        weight_mem[16'h0A5A] <= 0;
        weight_mem[16'h0A5B] <= 0;
        weight_mem[16'h0A5C] <= 0;
        weight_mem[16'h0A5D] <= 0;
        weight_mem[16'h0A5E] <= 0;
        weight_mem[16'h0A5F] <= 0;
        weight_mem[16'h0A60] <= 0;
        weight_mem[16'h0A61] <= 0;
        weight_mem[16'h0A62] <= 0;
        weight_mem[16'h0A63] <= 0;
        weight_mem[16'h0A64] <= 0;
        weight_mem[16'h0A65] <= 0;
        weight_mem[16'h0A66] <= 0;
        weight_mem[16'h0A67] <= 0;
        weight_mem[16'h0A68] <= 0;
        weight_mem[16'h0A69] <= 0;
        weight_mem[16'h0A6A] <= 0;
        weight_mem[16'h0A6B] <= 0;
        weight_mem[16'h0A6C] <= 0;
        weight_mem[16'h0A6D] <= 0;
        weight_mem[16'h0A6E] <= 0;
        weight_mem[16'h0A6F] <= 0;
        weight_mem[16'h0A70] <= 0;
        weight_mem[16'h0A71] <= 0;
        weight_mem[16'h0A72] <= 0;
        weight_mem[16'h0A73] <= 0;
        weight_mem[16'h0A74] <= 0;
        weight_mem[16'h0A75] <= 0;
        weight_mem[16'h0A76] <= 0;
        weight_mem[16'h0A77] <= 0;
        weight_mem[16'h0A78] <= 0;
        weight_mem[16'h0A79] <= 0;
        weight_mem[16'h0A7A] <= 0;
        weight_mem[16'h0A7B] <= 0;
        weight_mem[16'h0A7C] <= 0;
        weight_mem[16'h0A7D] <= 0;
        weight_mem[16'h0A7E] <= 0;
        weight_mem[16'h0A7F] <= 0;
        weight_mem[16'h0A80] <= 0;
        weight_mem[16'h0A81] <= 0;
        weight_mem[16'h0A82] <= 0;
        weight_mem[16'h0A83] <= 0;
        weight_mem[16'h0A84] <= 0;
        weight_mem[16'h0A85] <= 0;
        weight_mem[16'h0A86] <= 0;
        weight_mem[16'h0A87] <= 0;
        weight_mem[16'h0A88] <= 0;
        weight_mem[16'h0A89] <= 0;
        weight_mem[16'h0A8A] <= 0;
        weight_mem[16'h0A8B] <= 0;
        weight_mem[16'h0A8C] <= 0;
        weight_mem[16'h0A8D] <= 0;
        weight_mem[16'h0A8E] <= 0;
        weight_mem[16'h0A8F] <= 0;
        weight_mem[16'h0A90] <= 0;
        weight_mem[16'h0A91] <= 0;
        weight_mem[16'h0A92] <= 0;
        weight_mem[16'h0A93] <= 0;
        weight_mem[16'h0A94] <= 0;
        weight_mem[16'h0A95] <= 0;
        weight_mem[16'h0A96] <= 0;
        weight_mem[16'h0A97] <= 0;
        weight_mem[16'h0A98] <= 0;
        weight_mem[16'h0A99] <= 0;
        weight_mem[16'h0A9A] <= 0;
        weight_mem[16'h0A9B] <= 0;
        weight_mem[16'h0A9C] <= 0;
        weight_mem[16'h0A9D] <= 0;
        weight_mem[16'h0A9E] <= 0;
        weight_mem[16'h0A9F] <= 0;
        weight_mem[16'h0AA0] <= 0;
        weight_mem[16'h0AA1] <= 0;
        weight_mem[16'h0AA2] <= 0;
        weight_mem[16'h0AA3] <= 0;
        weight_mem[16'h0AA4] <= 0;
        weight_mem[16'h0AA5] <= 0;
        weight_mem[16'h0AA6] <= 0;
        weight_mem[16'h0AA7] <= 0;
        weight_mem[16'h0AA8] <= 0;
        weight_mem[16'h0AA9] <= 0;
        weight_mem[16'h0AAA] <= 0;
        weight_mem[16'h0AAB] <= 0;
        weight_mem[16'h0AAC] <= 0;
        weight_mem[16'h0AAD] <= 0;
        weight_mem[16'h0AAE] <= 0;
        weight_mem[16'h0AAF] <= 0;
        weight_mem[16'h0AB0] <= 0;
        weight_mem[16'h0AB1] <= 0;
        weight_mem[16'h0AB2] <= 0;
        weight_mem[16'h0AB3] <= 0;
        weight_mem[16'h0AB4] <= 0;
        weight_mem[16'h0AB5] <= 0;
        weight_mem[16'h0AB6] <= 0;
        weight_mem[16'h0AB7] <= 0;
        weight_mem[16'h0AB8] <= 0;
        weight_mem[16'h0AB9] <= 0;
        weight_mem[16'h0ABA] <= 0;
        weight_mem[16'h0ABB] <= 0;
        weight_mem[16'h0ABC] <= 0;
        weight_mem[16'h0ABD] <= 0;
        weight_mem[16'h0ABE] <= 0;
        weight_mem[16'h0ABF] <= 0;
        weight_mem[16'h0AC0] <= 0;
        weight_mem[16'h0AC1] <= 0;
        weight_mem[16'h0AC2] <= 0;
        weight_mem[16'h0AC3] <= 0;
        weight_mem[16'h0AC4] <= 0;
        weight_mem[16'h0AC5] <= 0;
        weight_mem[16'h0AC6] <= 0;
        weight_mem[16'h0AC7] <= 0;
        weight_mem[16'h0AC8] <= 0;
        weight_mem[16'h0AC9] <= 0;
        weight_mem[16'h0ACA] <= 0;
        weight_mem[16'h0ACB] <= 0;
        weight_mem[16'h0ACC] <= 0;
        weight_mem[16'h0ACD] <= 0;
        weight_mem[16'h0ACE] <= 0;
        weight_mem[16'h0ACF] <= 0;
        weight_mem[16'h0AD0] <= 0;
        weight_mem[16'h0AD1] <= 0;
        weight_mem[16'h0AD2] <= 0;
        weight_mem[16'h0AD3] <= 0;
        weight_mem[16'h0AD4] <= 0;
        weight_mem[16'h0AD5] <= 0;
        weight_mem[16'h0AD6] <= 0;
        weight_mem[16'h0AD7] <= 0;
        weight_mem[16'h0AD8] <= 0;
        weight_mem[16'h0AD9] <= 0;
        weight_mem[16'h0ADA] <= 0;
        weight_mem[16'h0ADB] <= 0;
        weight_mem[16'h0ADC] <= 0;
        weight_mem[16'h0ADD] <= 0;
        weight_mem[16'h0ADE] <= 0;
        weight_mem[16'h0ADF] <= 0;
        weight_mem[16'h0AE0] <= 0;
        weight_mem[16'h0AE1] <= 0;
        weight_mem[16'h0AE2] <= 0;
        weight_mem[16'h0AE3] <= 0;
        weight_mem[16'h0AE4] <= 0;
        weight_mem[16'h0AE5] <= 0;
        weight_mem[16'h0AE6] <= 0;
        weight_mem[16'h0AE7] <= 0;
        weight_mem[16'h0AE8] <= 0;
        weight_mem[16'h0AE9] <= 0;
        weight_mem[16'h0AEA] <= 0;
        weight_mem[16'h0AEB] <= 0;
        weight_mem[16'h0AEC] <= 0;
        weight_mem[16'h0AED] <= 0;
        weight_mem[16'h0AEE] <= 0;
        weight_mem[16'h0AEF] <= 0;
        weight_mem[16'h0AF0] <= 0;
        weight_mem[16'h0AF1] <= 0;
        weight_mem[16'h0AF2] <= 0;
        weight_mem[16'h0AF3] <= 0;
        weight_mem[16'h0AF4] <= 0;
        weight_mem[16'h0AF5] <= 0;
        weight_mem[16'h0AF6] <= 0;
        weight_mem[16'h0AF7] <= 0;
        weight_mem[16'h0AF8] <= 0;
        weight_mem[16'h0AF9] <= 0;
        weight_mem[16'h0AFA] <= 0;
        weight_mem[16'h0AFB] <= 0;
        weight_mem[16'h0AFC] <= 0;
        weight_mem[16'h0AFD] <= 0;
        weight_mem[16'h0AFE] <= 0;
        weight_mem[16'h0AFF] <= 0;
        weight_mem[16'h0B00] <= 0;
        weight_mem[16'h0B01] <= 0;
        weight_mem[16'h0B02] <= 0;
        weight_mem[16'h0B03] <= 0;
        weight_mem[16'h0B04] <= 0;
        weight_mem[16'h0B05] <= 0;
        weight_mem[16'h0B06] <= 0;
        weight_mem[16'h0B07] <= 0;
        weight_mem[16'h0B08] <= 0;
        weight_mem[16'h0B09] <= 0;
        weight_mem[16'h0B0A] <= 0;
        weight_mem[16'h0B0B] <= 0;
        weight_mem[16'h0B0C] <= 0;
        weight_mem[16'h0B0D] <= 0;
        weight_mem[16'h0B0E] <= 0;
        weight_mem[16'h0B0F] <= 0;
        weight_mem[16'h0B10] <= 0;
        weight_mem[16'h0B11] <= 0;
        weight_mem[16'h0B12] <= 0;
        weight_mem[16'h0B13] <= 0;
        weight_mem[16'h0B14] <= 0;
        weight_mem[16'h0B15] <= 0;
        weight_mem[16'h0B16] <= 0;
        weight_mem[16'h0B17] <= 0;
        weight_mem[16'h0B18] <= 0;
        weight_mem[16'h0B19] <= 0;
        weight_mem[16'h0B1A] <= 0;
        weight_mem[16'h0B1B] <= 0;
        weight_mem[16'h0B1C] <= 0;
        weight_mem[16'h0B1D] <= 0;
        weight_mem[16'h0B1E] <= 0;
        weight_mem[16'h0B1F] <= 0;
        weight_mem[16'h0B20] <= 0;
        weight_mem[16'h0B21] <= 0;
        weight_mem[16'h0B22] <= 0;
        weight_mem[16'h0B23] <= 0;
        weight_mem[16'h0B24] <= 0;
        weight_mem[16'h0B25] <= 0;
        weight_mem[16'h0B26] <= 0;
        weight_mem[16'h0B27] <= 0;
        weight_mem[16'h0B28] <= 0;
        weight_mem[16'h0B29] <= 0;
        weight_mem[16'h0B2A] <= 0;
        weight_mem[16'h0B2B] <= 0;
        weight_mem[16'h0B2C] <= 0;
        weight_mem[16'h0B2D] <= 0;
        weight_mem[16'h0B2E] <= 0;
        weight_mem[16'h0B2F] <= 0;
        weight_mem[16'h0B30] <= 0;
        weight_mem[16'h0B31] <= 0;
        weight_mem[16'h0B32] <= 0;
        weight_mem[16'h0B33] <= 0;
        weight_mem[16'h0B34] <= 0;
        weight_mem[16'h0B35] <= 0;
        weight_mem[16'h0B36] <= 0;
        weight_mem[16'h0B37] <= 0;
        weight_mem[16'h0B38] <= 0;
        weight_mem[16'h0B39] <= 0;
        weight_mem[16'h0B3A] <= 0;
        weight_mem[16'h0B3B] <= 0;
        weight_mem[16'h0B3C] <= 0;
        weight_mem[16'h0B3D] <= 0;
        weight_mem[16'h0B3E] <= 0;
        weight_mem[16'h0B3F] <= 0;
        weight_mem[16'h0B40] <= 0;
        weight_mem[16'h0B41] <= 0;
        weight_mem[16'h0B42] <= 0;
        weight_mem[16'h0B43] <= 0;
        weight_mem[16'h0B44] <= 0;
        weight_mem[16'h0B45] <= 0;
        weight_mem[16'h0B46] <= 0;
        weight_mem[16'h0B47] <= 0;
        weight_mem[16'h0B48] <= 0;
        weight_mem[16'h0B49] <= 0;
        weight_mem[16'h0B4A] <= 0;
        weight_mem[16'h0B4B] <= 0;
        weight_mem[16'h0B4C] <= 0;
        weight_mem[16'h0B4D] <= 0;
        weight_mem[16'h0B4E] <= 0;
        weight_mem[16'h0B4F] <= 0;
        weight_mem[16'h0B50] <= 0;
        weight_mem[16'h0B51] <= 0;
        weight_mem[16'h0B52] <= 0;
        weight_mem[16'h0B53] <= 0;
        weight_mem[16'h0B54] <= 0;
        weight_mem[16'h0B55] <= 0;
        weight_mem[16'h0B56] <= 0;
        weight_mem[16'h0B57] <= 0;
        weight_mem[16'h0B58] <= 0;
        weight_mem[16'h0B59] <= 0;
        weight_mem[16'h0B5A] <= 0;
        weight_mem[16'h0B5B] <= 0;
        weight_mem[16'h0B5C] <= 0;
        weight_mem[16'h0B5D] <= 0;
        weight_mem[16'h0B5E] <= 255;
        weight_mem[16'h0B5F] <= 0;
        weight_mem[16'h0B60] <= 0;
        weight_mem[16'h0B61] <= 0;
        weight_mem[16'h0B62] <= 0;
        weight_mem[16'h0B63] <= 0;
        weight_mem[16'h0B64] <= 0;
        weight_mem[16'h0B65] <= 0;
        weight_mem[16'h0B66] <= 0;
        weight_mem[16'h0B67] <= 0;
        weight_mem[16'h0B68] <= 0;
        weight_mem[16'h0B69] <= 0;
        weight_mem[16'h0B6A] <= 0;
        weight_mem[16'h0B6B] <= 0;
        weight_mem[16'h0B6C] <= 0;
        weight_mem[16'h0B6D] <= 0;
        weight_mem[16'h0B6E] <= 0;
        weight_mem[16'h0B6F] <= 0;
        weight_mem[16'h0B70] <= 0;
        weight_mem[16'h0B71] <= 0;
        weight_mem[16'h0B72] <= 0;
        weight_mem[16'h0B73] <= 253;
        weight_mem[16'h0B74] <= 0;
        weight_mem[16'h0B75] <= 1;
        weight_mem[16'h0B76] <= 0;
        weight_mem[16'h0B77] <= 0;
        weight_mem[16'h0B78] <= 0;
        weight_mem[16'h0B79] <= 0;
        weight_mem[16'h0B7A] <= 0;
        weight_mem[16'h0B7B] <= 0;
        weight_mem[16'h0B7C] <= 0;
        weight_mem[16'h0B7D] <= 0;
        weight_mem[16'h0B7E] <= 0;
        weight_mem[16'h0B7F] <= 0;
        weight_mem[16'h0B80] <= 0;
        weight_mem[16'h0B81] <= 0;
        weight_mem[16'h0B82] <= 0;
        weight_mem[16'h0B83] <= 0;
        weight_mem[16'h0B84] <= 0;
        weight_mem[16'h0B85] <= 0;
        weight_mem[16'h0B86] <= 0;
        weight_mem[16'h0B87] <= 0;
        weight_mem[16'h0B88] <= 0;
        weight_mem[16'h0B89] <= 0;
        weight_mem[16'h0B8A] <= 0;
        weight_mem[16'h0B8B] <= 0;
        weight_mem[16'h0B8C] <= 0;
        weight_mem[16'h0B8D] <= 0;
        weight_mem[16'h0B8E] <= 0;
        weight_mem[16'h0B8F] <= 0;
        weight_mem[16'h0B90] <= 0;
        weight_mem[16'h0B91] <= 0;
        weight_mem[16'h0B92] <= 0;
        weight_mem[16'h0B93] <= 0;
        weight_mem[16'h0B94] <= 0;
        weight_mem[16'h0B95] <= 0;
        weight_mem[16'h0B96] <= 0;
        weight_mem[16'h0B97] <= 0;
        weight_mem[16'h0B98] <= 0;
        weight_mem[16'h0B99] <= 0;
        weight_mem[16'h0B9A] <= 0;
        weight_mem[16'h0B9B] <= 0;
        weight_mem[16'h0B9C] <= 0;
        weight_mem[16'h0B9D] <= 0;
        weight_mem[16'h0B9E] <= 0;
        weight_mem[16'h0B9F] <= 0;
        weight_mem[16'h0BA0] <= 0;
        weight_mem[16'h0BA1] <= 0;
        weight_mem[16'h0BA2] <= 0;
        weight_mem[16'h0BA3] <= 0;
        weight_mem[16'h0BA4] <= 0;
        weight_mem[16'h0BA5] <= 0;
        weight_mem[16'h0BA6] <= 0;
        weight_mem[16'h0BA7] <= 0;
        weight_mem[16'h0BA8] <= 0;
        weight_mem[16'h0BA9] <= 0;
        weight_mem[16'h0BAA] <= 0;
        weight_mem[16'h0BAB] <= 0;
        weight_mem[16'h0BAC] <= 0;
        weight_mem[16'h0BAD] <= 0;
        weight_mem[16'h0BAE] <= 0;
        weight_mem[16'h0BAF] <= 0;

        // layer 1 neuron 6
        weight_mem[16'h0C00] <= 243;
        weight_mem[16'h0C01] <= 14;
        weight_mem[16'h0C02] <= 1;
        weight_mem[16'h0C03] <= 7;
        weight_mem[16'h0C04] <= 5;
        weight_mem[16'h0C05] <= 242;
        weight_mem[16'h0C06] <= 244;
        weight_mem[16'h0C07] <= 249;
        weight_mem[16'h0C08] <= 10;
        weight_mem[16'h0C09] <= 243;
        weight_mem[16'h0C0A] <= 255;
        weight_mem[16'h0C0B] <= 253;
        weight_mem[16'h0C0C] <= 0;
        weight_mem[16'h0C0D] <= 10;
        weight_mem[16'h0C0E] <= 255;
        weight_mem[16'h0C0F] <= 13;
        weight_mem[16'h0C10] <= 15;
        weight_mem[16'h0C11] <= 253;
        weight_mem[16'h0C12] <= 241;
        weight_mem[16'h0C13] <= 2;
        weight_mem[16'h0C14] <= 244;
        weight_mem[16'h0C15] <= 253;
        weight_mem[16'h0C16] <= 254;
        weight_mem[16'h0C17] <= 241;
        weight_mem[16'h0C18] <= 9;
        weight_mem[16'h0C19] <= 5;
        weight_mem[16'h0C1A] <= 8;
        weight_mem[16'h0C1B] <= 15;
        weight_mem[16'h0C1C] <= 246;
        weight_mem[16'h0C1D] <= 4;
        weight_mem[16'h0C1E] <= 245;
        weight_mem[16'h0C1F] <= 10;
        weight_mem[16'h0C20] <= 14;
        weight_mem[16'h0C21] <= 19;
        weight_mem[16'h0C22] <= 5;
        weight_mem[16'h0C23] <= 21;
        weight_mem[16'h0C24] <= 26;
        weight_mem[16'h0C25] <= 11;
        weight_mem[16'h0C26] <= 2;
        weight_mem[16'h0C27] <= 0;
        weight_mem[16'h0C28] <= 4;
        weight_mem[16'h0C29] <= 20;
        weight_mem[16'h0C2A] <= 9;
        weight_mem[16'h0C2B] <= 15;
        weight_mem[16'h0C2C] <= 245;
        weight_mem[16'h0C2D] <= 8;
        weight_mem[16'h0C2E] <= 244;
        weight_mem[16'h0C2F] <= 8;
        weight_mem[16'h0C30] <= 246;
        weight_mem[16'h0C31] <= 250;
        weight_mem[16'h0C32] <= 250;
        weight_mem[16'h0C33] <= 2;
        weight_mem[16'h0C34] <= 3;
        weight_mem[16'h0C35] <= 12;
        weight_mem[16'h0C36] <= 252;
        weight_mem[16'h0C37] <= 18;
        weight_mem[16'h0C38] <= 26;
        weight_mem[16'h0C39] <= 37;
        weight_mem[16'h0C3A] <= 31;
        weight_mem[16'h0C3B] <= 23;
        weight_mem[16'h0C3C] <= 34;
        weight_mem[16'h0C3D] <= 24;
        weight_mem[16'h0C3E] <= 10;
        weight_mem[16'h0C3F] <= 21;
        weight_mem[16'h0C40] <= 23;
        weight_mem[16'h0C41] <= 15;
        weight_mem[16'h0C42] <= 13;
        weight_mem[16'h0C43] <= 22;
        weight_mem[16'h0C44] <= 18;
        weight_mem[16'h0C45] <= 14;
        weight_mem[16'h0C46] <= 247;
        weight_mem[16'h0C47] <= 251;
        weight_mem[16'h0C48] <= 10;
        weight_mem[16'h0C49] <= 10;
        weight_mem[16'h0C4A] <= 252;
        weight_mem[16'h0C4B] <= 13;
        weight_mem[16'h0C4C] <= 16;
        weight_mem[16'h0C4D] <= 10;
        weight_mem[16'h0C4E] <= 19;
        weight_mem[16'h0C4F] <= 54;
        weight_mem[16'h0C50] <= 39;
        weight_mem[16'h0C51] <= 57;
        weight_mem[16'h0C52] <= 86;
        weight_mem[16'h0C53] <= 73;
        weight_mem[16'h0C54] <= 72;
        weight_mem[16'h0C55] <= 78;
        weight_mem[16'h0C56] <= 98;
        weight_mem[16'h0C57] <= 75;
        weight_mem[16'h0C58] <= 79;
        weight_mem[16'h0C59] <= 52;
        weight_mem[16'h0C5A] <= 23;
        weight_mem[16'h0C5B] <= 255;
        weight_mem[16'h0C5C] <= 255;
        weight_mem[16'h0C5D] <= 254;
        weight_mem[16'h0C5E] <= 252;
        weight_mem[16'h0C5F] <= 1;
        weight_mem[16'h0C60] <= 241;
        weight_mem[16'h0C61] <= 15;
        weight_mem[16'h0C62] <= 0;
        weight_mem[16'h0C63] <= 4;
        weight_mem[16'h0C64] <= 4;
        weight_mem[16'h0C65] <= 255;
        weight_mem[16'h0C66] <= 255;
        weight_mem[16'h0C67] <= 3;
        weight_mem[16'h0C68] <= 248;
        weight_mem[16'h0C69] <= 5;
        weight_mem[16'h0C6A] <= 252;
        weight_mem[16'h0C6B] <= 18;
        weight_mem[16'h0C6C] <= 26;
        weight_mem[16'h0C6D] <= 39;
        weight_mem[16'h0C6E] <= 22;
        weight_mem[16'h0C6F] <= 251;
        weight_mem[16'h0C70] <= 252;
        weight_mem[16'h0C71] <= 235;
        weight_mem[16'h0C72] <= 236;
        weight_mem[16'h0C73] <= 198;
        weight_mem[16'h0C74] <= 205;
        weight_mem[16'h0C75] <= 241;
        weight_mem[16'h0C76] <= 231;
        weight_mem[16'h0C77] <= 0;
        weight_mem[16'h0C78] <= 252;
        weight_mem[16'h0C79] <= 238;
        weight_mem[16'h0C7A] <= 4;
        weight_mem[16'h0C7B] <= 255;
        weight_mem[16'h0C7C] <= 249;
        weight_mem[16'h0C7D] <= 238;
        weight_mem[16'h0C7E] <= 228;
        weight_mem[16'h0C7F] <= 213;
        weight_mem[16'h0C80] <= 214;
        weight_mem[16'h0C81] <= 224;
        weight_mem[16'h0C82] <= 187;
        weight_mem[16'h0C83] <= 179;
        weight_mem[16'h0C84] <= 202;
        weight_mem[16'h0C85] <= 196;
        weight_mem[16'h0C86] <= 194;
        weight_mem[16'h0C87] <= 207;
        weight_mem[16'h0C88] <= 214;
        weight_mem[16'h0C89] <= 184;
        weight_mem[16'h0C8A] <= 175;
        weight_mem[16'h0C8B] <= 162;
        weight_mem[16'h0C8C] <= 148;
        weight_mem[16'h0C8D] <= 191;
        weight_mem[16'h0C8E] <= 225;
        weight_mem[16'h0C8F] <= 249;
        weight_mem[16'h0C90] <= 248;
        weight_mem[16'h0C91] <= 243;
        weight_mem[16'h0C92] <= 226;
        weight_mem[16'h0C93] <= 225;
        weight_mem[16'h0C94] <= 229;
        weight_mem[16'h0C95] <= 227;
        weight_mem[16'h0C96] <= 245;
        weight_mem[16'h0C97] <= 242;
        weight_mem[16'h0C98] <= 232;
        weight_mem[16'h0C99] <= 205;
        weight_mem[16'h0C9A] <= 171;
        weight_mem[16'h0C9B] <= 128;
        weight_mem[16'h0C9C] <= 139;
        weight_mem[16'h0C9D] <= 168;
        weight_mem[16'h0C9E] <= 206;
        weight_mem[16'h0C9F] <= 212;
        weight_mem[16'h0CA0] <= 228;
        weight_mem[16'h0CA1] <= 177;
        weight_mem[16'h0CA2] <= 180;
        weight_mem[16'h0CA3] <= 172;
        weight_mem[16'h0CA4] <= 175;
        weight_mem[16'h0CA5] <= 182;
        weight_mem[16'h0CA6] <= 221;
        weight_mem[16'h0CA7] <= 5;
        weight_mem[16'h0CA8] <= 250;
        weight_mem[16'h0CA9] <= 238;
        weight_mem[16'h0CAA] <= 1;
        weight_mem[16'h0CAB] <= 226;
        weight_mem[16'h0CAC] <= 230;
        weight_mem[16'h0CAD] <= 243;
        weight_mem[16'h0CAE] <= 242;
        weight_mem[16'h0CAF] <= 237;
        weight_mem[16'h0CB0] <= 239;
        weight_mem[16'h0CB1] <= 203;
        weight_mem[16'h0CB2] <= 167;
        weight_mem[16'h0CB3] <= 132;
        weight_mem[16'h0CB4] <= 179;
        weight_mem[16'h0CB5] <= 206;
        weight_mem[16'h0CB6] <= 236;
        weight_mem[16'h0CB7] <= 243;
        weight_mem[16'h0CB8] <= 13;
        weight_mem[16'h0CB9] <= 253;
        weight_mem[16'h0CBA] <= 237;
        weight_mem[16'h0CBB] <= 3;
        weight_mem[16'h0CBC] <= 233;
        weight_mem[16'h0CBD] <= 229;
        weight_mem[16'h0CBE] <= 245;
        weight_mem[16'h0CBF] <= 250;
        weight_mem[16'h0CC0] <= 242;
        weight_mem[16'h0CC1] <= 3;
        weight_mem[16'h0CC2] <= 232;
        weight_mem[16'h0CC3] <= 0;
        weight_mem[16'h0CC4] <= 232;
        weight_mem[16'h0CC5] <= 247;
        weight_mem[16'h0CC6] <= 232;
        weight_mem[16'h0CC7] <= 234;
        weight_mem[16'h0CC8] <= 0;
        weight_mem[16'h0CC9] <= 10;
        weight_mem[16'h0CCA] <= 18;
        weight_mem[16'h0CCB] <= 40;
        weight_mem[16'h0CCC] <= 15;
        weight_mem[16'h0CCD] <= 49;
        weight_mem[16'h0CCE] <= 44;
        weight_mem[16'h0CCF] <= 48;
        weight_mem[16'h0CD0] <= 47;
        weight_mem[16'h0CD1] <= 16;
        weight_mem[16'h0CD2] <= 24;
        weight_mem[16'h0CD3] <= 22;
        weight_mem[16'h0CD4] <= 20;
        weight_mem[16'h0CD5] <= 249;
        weight_mem[16'h0CD6] <= 240;
        weight_mem[16'h0CD7] <= 244;
        weight_mem[16'h0CD8] <= 13;
        weight_mem[16'h0CD9] <= 242;
        weight_mem[16'h0CDA] <= 255;
        weight_mem[16'h0CDB] <= 11;
        weight_mem[16'h0CDC] <= 8;
        weight_mem[16'h0CDD] <= 4;
        weight_mem[16'h0CDE] <= 0;
        weight_mem[16'h0CDF] <= 8;
        weight_mem[16'h0CE0] <= 248;
        weight_mem[16'h0CE1] <= 18;
        weight_mem[16'h0CE2] <= 40;
        weight_mem[16'h0CE3] <= 71;
        weight_mem[16'h0CE4] <= 54;
        weight_mem[16'h0CE5] <= 29;
        weight_mem[16'h0CE6] <= 31;
        weight_mem[16'h0CE7] <= 17;
        weight_mem[16'h0CE8] <= 5;
        weight_mem[16'h0CE9] <= 241;
        weight_mem[16'h0CEA] <= 0;
        weight_mem[16'h0CEB] <= 4;
        weight_mem[16'h0CEC] <= 13;
        weight_mem[16'h0CED] <= 247;
        weight_mem[16'h0CEE] <= 242;
        weight_mem[16'h0CEF] <= 9;
        weight_mem[16'h0CF0] <= 4;
        weight_mem[16'h0CF1] <= 253;
        weight_mem[16'h0CF2] <= 251;
        weight_mem[16'h0CF3] <= 12;
        weight_mem[16'h0CF4] <= 3;
        weight_mem[16'h0CF5] <= 22;
        weight_mem[16'h0CF6] <= 21;
        weight_mem[16'h0CF7] <= 17;
        weight_mem[16'h0CF8] <= 10;
        weight_mem[16'h0CF9] <= 46;
        weight_mem[16'h0CFA] <= 26;
        weight_mem[16'h0CFB] <= 50;
        weight_mem[16'h0CFC] <= 50;
        weight_mem[16'h0CFD] <= 253;
        weight_mem[16'h0CFE] <= 244;
        weight_mem[16'h0CFF] <= 218;
        weight_mem[16'h0D00] <= 236;
        weight_mem[16'h0D01] <= 251;
        weight_mem[16'h0D02] <= 0;
        weight_mem[16'h0D03] <= 1;
        weight_mem[16'h0D04] <= 17;
        weight_mem[16'h0D05] <= 14;
        weight_mem[16'h0D06] <= 16;
        weight_mem[16'h0D07] <= 248;
        weight_mem[16'h0D08] <= 11;
        weight_mem[16'h0D09] <= 15;
        weight_mem[16'h0D0A] <= 13;
        weight_mem[16'h0D0B] <= 14;
        weight_mem[16'h0D0C] <= 1;
        weight_mem[16'h0D0D] <= 243;
        weight_mem[16'h0D0E] <= 10;
        weight_mem[16'h0D0F] <= 36;
        weight_mem[16'h0D10] <= 42;
        weight_mem[16'h0D11] <= 62;
        weight_mem[16'h0D12] <= 58;
        weight_mem[16'h0D13] <= 23;
        weight_mem[16'h0D14] <= 237;
        weight_mem[16'h0D15] <= 219;
        weight_mem[16'h0D16] <= 240;
        weight_mem[16'h0D17] <= 15;
        weight_mem[16'h0D18] <= 41;
        weight_mem[16'h0D19] <= 24;
        weight_mem[16'h0D1A] <= 27;
        weight_mem[16'h0D1B] <= 41;
        weight_mem[16'h0D1C] <= 39;
        weight_mem[16'h0D1D] <= 27;
        weight_mem[16'h0D1E] <= 12;
        weight_mem[16'h0D1F] <= 244;
        weight_mem[16'h0D20] <= 5;
        weight_mem[16'h0D21] <= 246;
        weight_mem[16'h0D22] <= 15;
        weight_mem[16'h0D23] <= 3;
        weight_mem[16'h0D24] <= 5;
        weight_mem[16'h0D25] <= 235;
        weight_mem[16'h0D26] <= 249;
        weight_mem[16'h0D27] <= 22;
        weight_mem[16'h0D28] <= 41;
        weight_mem[16'h0D29] <= 67;
        weight_mem[16'h0D2A] <= 45;
        weight_mem[16'h0D2B] <= 236;
        weight_mem[16'h0D2C] <= 231;
        weight_mem[16'h0D2D] <= 29;
        weight_mem[16'h0D2E] <= 52;
        weight_mem[16'h0D2F] <= 66;
        weight_mem[16'h0D30] <= 42;
        weight_mem[16'h0D31] <= 52;
        weight_mem[16'h0D32] <= 74;
        weight_mem[16'h0D33] <= 62;
        weight_mem[16'h0D34] <= 43;
        weight_mem[16'h0D35] <= 6;
        weight_mem[16'h0D36] <= 244;
        weight_mem[16'h0D37] <= 245;
        weight_mem[16'h0D38] <= 0;
        weight_mem[16'h0D39] <= 8;
        weight_mem[16'h0D3A] <= 243;
        weight_mem[16'h0D3B] <= 12;
        weight_mem[16'h0D3C] <= 8;
        weight_mem[16'h0D3D] <= 13;
        weight_mem[16'h0D3E] <= 18;
        weight_mem[16'h0D3F] <= 24;
        weight_mem[16'h0D40] <= 55;
        weight_mem[16'h0D41] <= 62;
        weight_mem[16'h0D42] <= 23;
        weight_mem[16'h0D43] <= 1;
        weight_mem[16'h0D44] <= 31;
        weight_mem[16'h0D45] <= 42;
        weight_mem[16'h0D46] <= 63;
        weight_mem[16'h0D47] <= 66;
        weight_mem[16'h0D48] <= 68;
        weight_mem[16'h0D49] <= 81;
        weight_mem[16'h0D4A] <= 50;
        weight_mem[16'h0D4B] <= 35;
        weight_mem[16'h0D4C] <= 25;
        weight_mem[16'h0D4D] <= 246;
        weight_mem[16'h0D4E] <= 243;
        weight_mem[16'h0D4F] <= 252;
        weight_mem[16'h0D50] <= 2;
        weight_mem[16'h0D51] <= 4;
        weight_mem[16'h0D52] <= 255;
        weight_mem[16'h0D53] <= 249;
        weight_mem[16'h0D54] <= 11;
        weight_mem[16'h0D55] <= 2;
        weight_mem[16'h0D56] <= 14;
        weight_mem[16'h0D57] <= 22;
        weight_mem[16'h0D58] <= 25;
        weight_mem[16'h0D59] <= 44;
        weight_mem[16'h0D5A] <= 39;
        weight_mem[16'h0D5B] <= 57;
        weight_mem[16'h0D5C] <= 35;
        weight_mem[16'h0D5D] <= 44;
        weight_mem[16'h0D5E] <= 58;
        weight_mem[16'h0D5F] <= 61;
        weight_mem[16'h0D60] <= 74;
        weight_mem[16'h0D61] <= 78;
        weight_mem[16'h0D62] <= 39;
        weight_mem[16'h0D63] <= 26;
        weight_mem[16'h0D64] <= 250;
        weight_mem[16'h0D65] <= 14;
        weight_mem[16'h0D66] <= 251;
        weight_mem[16'h0D67] <= 0;
        weight_mem[16'h0D68] <= 250;
        weight_mem[16'h0D69] <= 254;
        weight_mem[16'h0D6A] <= 1;
        weight_mem[16'h0D6B] <= 12;
        weight_mem[16'h0D6C] <= 250;
        weight_mem[16'h0D6D] <= 238;
        weight_mem[16'h0D6E] <= 239;
        weight_mem[16'h0D6F] <= 245;
        weight_mem[16'h0D70] <= 234;
        weight_mem[16'h0D71] <= 222;
        weight_mem[16'h0D72] <= 222;
        weight_mem[16'h0D73] <= 252;
        weight_mem[16'h0D74] <= 234;
        weight_mem[16'h0D75] <= 255;
        weight_mem[16'h0D76] <= 12;
        weight_mem[16'h0D77] <= 8;
        weight_mem[16'h0D78] <= 17;
        weight_mem[16'h0D79] <= 22;
        weight_mem[16'h0D7A] <= 28;
        weight_mem[16'h0D7B] <= 13;
        weight_mem[16'h0D7C] <= 10;
        weight_mem[16'h0D7D] <= 6;
        weight_mem[16'h0D7E] <= 242;
        weight_mem[16'h0D7F] <= 249;
        weight_mem[16'h0D80] <= 252;
        weight_mem[16'h0D81] <= 9;
        weight_mem[16'h0D82] <= 247;
        weight_mem[16'h0D83] <= 237;
        weight_mem[16'h0D84] <= 244;
        weight_mem[16'h0D85] <= 238;
        weight_mem[16'h0D86] <= 227;
        weight_mem[16'h0D87] <= 204;
        weight_mem[16'h0D88] <= 221;
        weight_mem[16'h0D89] <= 214;
        weight_mem[16'h0D8A] <= 199;
        weight_mem[16'h0D8B] <= 186;
        weight_mem[16'h0D8C] <= 195;
        weight_mem[16'h0D8D] <= 189;
        weight_mem[16'h0D8E] <= 206;
        weight_mem[16'h0D8F] <= 232;
        weight_mem[16'h0D90] <= 248;
        weight_mem[16'h0D91] <= 14;
        weight_mem[16'h0D92] <= 255;
        weight_mem[16'h0D93] <= 11;
        weight_mem[16'h0D94] <= 255;
        weight_mem[16'h0D95] <= 3;
        weight_mem[16'h0D96] <= 241;
        weight_mem[16'h0D97] <= 13;
        weight_mem[16'h0D98] <= 6;
        weight_mem[16'h0D99] <= 15;
        weight_mem[16'h0D9A] <= 240;
        weight_mem[16'h0D9B] <= 246;
        weight_mem[16'h0D9C] <= 9;
        weight_mem[16'h0D9D] <= 10;
        weight_mem[16'h0D9E] <= 246;
        weight_mem[16'h0D9F] <= 1;
        weight_mem[16'h0DA0] <= 232;
        weight_mem[16'h0DA1] <= 231;
        weight_mem[16'h0DA2] <= 233;
        weight_mem[16'h0DA3] <= 241;
        weight_mem[16'h0DA4] <= 249;
        weight_mem[16'h0DA5] <= 249;
        weight_mem[16'h0DA6] <= 0;
        weight_mem[16'h0DA7] <= 252;
        weight_mem[16'h0DA8] <= 244;
        weight_mem[16'h0DA9] <= 246;
        weight_mem[16'h0DAA] <= 252;
        weight_mem[16'h0DAB] <= 1;
        weight_mem[16'h0DAC] <= 241;
        weight_mem[16'h0DAD] <= 12;
        weight_mem[16'h0DAE] <= 249;
        weight_mem[16'h0DAF] <= 2;

        // layer 1 neuron 7
        weight_mem[16'h0E00] <= 180;
        weight_mem[16'h0E01] <= 180;
        weight_mem[16'h0E02] <= 180;
        weight_mem[16'h0E03] <= 180;
        weight_mem[16'h0E04] <= 180;
        weight_mem[16'h0E05] <= 180;
        weight_mem[16'h0E06] <= 180;
        weight_mem[16'h0E07] <= 180;
        weight_mem[16'h0E08] <= 180;
        weight_mem[16'h0E09] <= 180;
        weight_mem[16'h0E0A] <= 180;
        weight_mem[16'h0E0B] <= 180;
        weight_mem[16'h0E0C] <= 178;
        weight_mem[16'h0E0D] <= 177;
        weight_mem[16'h0E0E] <= 179;
        weight_mem[16'h0E0F] <= 180;
        weight_mem[16'h0E10] <= 180;
        weight_mem[16'h0E11] <= 180;
        weight_mem[16'h0E12] <= 180;
        weight_mem[16'h0E13] <= 180;
        weight_mem[16'h0E14] <= 180;
        weight_mem[16'h0E15] <= 180;
        weight_mem[16'h0E16] <= 180;
        weight_mem[16'h0E17] <= 180;
        weight_mem[16'h0E18] <= 180;
        weight_mem[16'h0E19] <= 180;
        weight_mem[16'h0E1A] <= 180;
        weight_mem[16'h0E1B] <= 180;
        weight_mem[16'h0E1C] <= 180;
        weight_mem[16'h0E1D] <= 180;
        weight_mem[16'h0E1E] <= 180;
        weight_mem[16'h0E1F] <= 180;
        weight_mem[16'h0E20] <= 179;
        weight_mem[16'h0E21] <= 179;
        weight_mem[16'h0E22] <= 179;
        weight_mem[16'h0E23] <= 178;
        weight_mem[16'h0E24] <= 174;
        weight_mem[16'h0E25] <= 172;
        weight_mem[16'h0E26] <= 174;
        weight_mem[16'h0E27] <= 177;
        weight_mem[16'h0E28] <= 178;
        weight_mem[16'h0E29] <= 179;
        weight_mem[16'h0E2A] <= 180;
        weight_mem[16'h0E2B] <= 180;
        weight_mem[16'h0E2C] <= 181;
        weight_mem[16'h0E2D] <= 180;
        weight_mem[16'h0E2E] <= 180;
        weight_mem[16'h0E2F] <= 180;
        weight_mem[16'h0E30] <= 180;
        weight_mem[16'h0E31] <= 180;
        weight_mem[16'h0E32] <= 180;
        weight_mem[16'h0E33] <= 180;
        weight_mem[16'h0E34] <= 180;
        weight_mem[16'h0E35] <= 180;
        weight_mem[16'h0E36] <= 180;
        weight_mem[16'h0E37] <= 179;
        weight_mem[16'h0E38] <= 176;
        weight_mem[16'h0E39] <= 172;
        weight_mem[16'h0E3A] <= 168;
        weight_mem[16'h0E3B] <= 165;
        weight_mem[16'h0E3C] <= 165;
        weight_mem[16'h0E3D] <= 162;
        weight_mem[16'h0E3E] <= 157;
        weight_mem[16'h0E3F] <= 165;
        weight_mem[16'h0E40] <= 172;
        weight_mem[16'h0E41] <= 178;
        weight_mem[16'h0E42] <= 182;
        weight_mem[16'h0E43] <= 184;
        weight_mem[16'h0E44] <= 190;
        weight_mem[16'h0E45] <= 185;
        weight_mem[16'h0E46] <= 180;
        weight_mem[16'h0E47] <= 180;
        weight_mem[16'h0E48] <= 180;
        weight_mem[16'h0E49] <= 180;
        weight_mem[16'h0E4A] <= 180;
        weight_mem[16'h0E4B] <= 180;
        weight_mem[16'h0E4C] <= 179;
        weight_mem[16'h0E4D] <= 179;
        weight_mem[16'h0E4E] <= 180;
        weight_mem[16'h0E4F] <= 172;
        weight_mem[16'h0E50] <= 160;
        weight_mem[16'h0E51] <= 151;
        weight_mem[16'h0E52] <= 152;
        weight_mem[16'h0E53] <= 151;
        weight_mem[16'h0E54] <= 140;
        weight_mem[16'h0E55] <= 129;
        weight_mem[16'h0E56] <= 132;
        weight_mem[16'h0E57] <= 157;
        weight_mem[16'h0E58] <= 180;
        weight_mem[16'h0E59] <= 185;
        weight_mem[16'h0E5A] <= 189;
        weight_mem[16'h0E5B] <= 186;
        weight_mem[16'h0E5C] <= 185;
        weight_mem[16'h0E5D] <= 182;
        weight_mem[16'h0E5E] <= 180;
        weight_mem[16'h0E5F] <= 180;
        weight_mem[16'h0E60] <= 180;
        weight_mem[16'h0E61] <= 180;
        weight_mem[16'h0E62] <= 180;
        weight_mem[16'h0E63] <= 180;
        weight_mem[16'h0E64] <= 182;
        weight_mem[16'h0E65] <= 190;
        weight_mem[16'h0E66] <= 188;
        weight_mem[16'h0E67] <= 175;
        weight_mem[16'h0E68] <= 164;
        weight_mem[16'h0E69] <= 164;
        weight_mem[16'h0E6A] <= 181;
        weight_mem[16'h0E6B] <= 187;
        weight_mem[16'h0E6C] <= 183;
        weight_mem[16'h0E6D] <= 171;
        weight_mem[16'h0E6E] <= 165;
        weight_mem[16'h0E6F] <= 170;
        weight_mem[16'h0E70] <= 174;
        weight_mem[16'h0E71] <= 171;
        weight_mem[16'h0E72] <= 182;
        weight_mem[16'h0E73] <= 181;
        weight_mem[16'h0E74] <= 175;
        weight_mem[16'h0E75] <= 175;
        weight_mem[16'h0E76] <= 179;
        weight_mem[16'h0E77] <= 180;
        weight_mem[16'h0E78] <= 180;
        weight_mem[16'h0E79] <= 180;
        weight_mem[16'h0E7A] <= 181;
        weight_mem[16'h0E7B] <= 183;
        weight_mem[16'h0E7C] <= 188;
        weight_mem[16'h0E7D] <= 194;
        weight_mem[16'h0E7E] <= 183;
        weight_mem[16'h0E7F] <= 183;
        weight_mem[16'h0E80] <= 188;
        weight_mem[16'h0E81] <= 176;
        weight_mem[16'h0E82] <= 188;
        weight_mem[16'h0E83] <= 208;
        weight_mem[16'h0E84] <= 223;
        weight_mem[16'h0E85] <= 214;
        weight_mem[16'h0E86] <= 194;
        weight_mem[16'h0E87] <= 184;
        weight_mem[16'h0E88] <= 148;
        weight_mem[16'h0E89] <= 138;
        weight_mem[16'h0E8A] <= 168;
        weight_mem[16'h0E8B] <= 176;
        weight_mem[16'h0E8C] <= 176;
        weight_mem[16'h0E8D] <= 176;
        weight_mem[16'h0E8E] <= 179;
        weight_mem[16'h0E8F] <= 180;
        weight_mem[16'h0E90] <= 180;
        weight_mem[16'h0E91] <= 180;
        weight_mem[16'h0E92] <= 180;
        weight_mem[16'h0E93] <= 181;
        weight_mem[16'h0E94] <= 182;
        weight_mem[16'h0E95] <= 178;
        weight_mem[16'h0E96] <= 175;
        weight_mem[16'h0E97] <= 186;
        weight_mem[16'h0E98] <= 184;
        weight_mem[16'h0E99] <= 174;
        weight_mem[16'h0E9A] <= 177;
        weight_mem[16'h0E9B] <= 203;
        weight_mem[16'h0E9C] <= 220;
        weight_mem[16'h0E9D] <= 214;
        weight_mem[16'h0E9E] <= 193;
        weight_mem[16'h0E9F] <= 171;
        weight_mem[16'h0EA0] <= 150;
        weight_mem[16'h0EA1] <= 151;
        weight_mem[16'h0EA2] <= 174;
        weight_mem[16'h0EA3] <= 175;
        weight_mem[16'h0EA4] <= 176;
        weight_mem[16'h0EA5] <= 176;
        weight_mem[16'h0EA6] <= 178;
        weight_mem[16'h0EA7] <= 180;
        weight_mem[16'h0EA8] <= 180;
        weight_mem[16'h0EA9] <= 180;
        weight_mem[16'h0EAA] <= 179;
        weight_mem[16'h0EAB] <= 178;
        weight_mem[16'h0EAC] <= 176;
        weight_mem[16'h0EAD] <= 175;
        weight_mem[16'h0EAE] <= 179;
        weight_mem[16'h0EAF] <= 181;
        weight_mem[16'h0EB0] <= 188;
        weight_mem[16'h0EB1] <= 192;
        weight_mem[16'h0EB2] <= 191;
        weight_mem[16'h0EB3] <= 200;
        weight_mem[16'h0EB4] <= 195;
        weight_mem[16'h0EB5] <= 184;
        weight_mem[16'h0EB6] <= 174;
        weight_mem[16'h0EB7] <= 157;
        weight_mem[16'h0EB8] <= 156;
        weight_mem[16'h0EB9] <= 170;
        weight_mem[16'h0EBA] <= 174;
        weight_mem[16'h0EBB] <= 174;
        weight_mem[16'h0EBC] <= 178;
        weight_mem[16'h0EBD] <= 179;
        weight_mem[16'h0EBE] <= 179;
        weight_mem[16'h0EBF] <= 179;
        weight_mem[16'h0EC0] <= 180;
        weight_mem[16'h0EC1] <= 180;
        weight_mem[16'h0EC2] <= 179;
        weight_mem[16'h0EC3] <= 178;
        weight_mem[16'h0EC4] <= 177;
        weight_mem[16'h0EC5] <= 172;
        weight_mem[16'h0EC6] <= 175;
        weight_mem[16'h0EC7] <= 183;
        weight_mem[16'h0EC8] <= 190;
        weight_mem[16'h0EC9] <= 197;
        weight_mem[16'h0ECA] <= 198;
        weight_mem[16'h0ECB] <= 198;
        weight_mem[16'h0ECC] <= 193;
        weight_mem[16'h0ECD] <= 186;
        weight_mem[16'h0ECE] <= 174;
        weight_mem[16'h0ECF] <= 151;
        weight_mem[16'h0ED0] <= 136;
        weight_mem[16'h0ED1] <= 161;
        weight_mem[16'h0ED2] <= 164;
        weight_mem[16'h0ED3] <= 165;
        weight_mem[16'h0ED4] <= 175;
        weight_mem[16'h0ED5] <= 179;
        weight_mem[16'h0ED6] <= 180;
        weight_mem[16'h0ED7] <= 180;
        weight_mem[16'h0ED8] <= 180;
        weight_mem[16'h0ED9] <= 180;
        weight_mem[16'h0EDA] <= 180;
        weight_mem[16'h0EDB] <= 179;
        weight_mem[16'h0EDC] <= 175;
        weight_mem[16'h0EDD] <= 162;
        weight_mem[16'h0EDE] <= 169;
        weight_mem[16'h0EDF] <= 181;
        weight_mem[16'h0EE0] <= 182;
        weight_mem[16'h0EE1] <= 181;
        weight_mem[16'h0EE2] <= 185;
        weight_mem[16'h0EE3] <= 198;
        weight_mem[16'h0EE4] <= 201;
        weight_mem[16'h0EE5] <= 186;
        weight_mem[16'h0EE6] <= 176;
        weight_mem[16'h0EE7] <= 152;
        weight_mem[16'h0EE8] <= 129;
        weight_mem[16'h0EE9] <= 150;
        weight_mem[16'h0EEA] <= 166;
        weight_mem[16'h0EEB] <= 170;
        weight_mem[16'h0EEC] <= 178;
        weight_mem[16'h0EED] <= 180;
        weight_mem[16'h0EEE] <= 180;
        weight_mem[16'h0EEF] <= 180;
        weight_mem[16'h0EF0] <= 180;
        weight_mem[16'h0EF1] <= 180;
        weight_mem[16'h0EF2] <= 180;
        weight_mem[16'h0EF3] <= 176;
        weight_mem[16'h0EF4] <= 165;
        weight_mem[16'h0EF5] <= 153;
        weight_mem[16'h0EF6] <= 156;
        weight_mem[16'h0EF7] <= 157;
        weight_mem[16'h0EF8] <= 155;
        weight_mem[16'h0EF9] <= 158;
        weight_mem[16'h0EFA] <= 173;
        weight_mem[16'h0EFB] <= 182;
        weight_mem[16'h0EFC] <= 200;
        weight_mem[16'h0EFD] <= 209;
        weight_mem[16'h0EFE] <= 191;
        weight_mem[16'h0EFF] <= 158;
        weight_mem[16'h0F00] <= 133;
        weight_mem[16'h0F01] <= 145;
        weight_mem[16'h0F02] <= 169;
        weight_mem[16'h0F03] <= 187;
        weight_mem[16'h0F04] <= 186;
        weight_mem[16'h0F05] <= 181;
        weight_mem[16'h0F06] <= 180;
        weight_mem[16'h0F07] <= 180;
        weight_mem[16'h0F08] <= 180;
        weight_mem[16'h0F09] <= 180;
        weight_mem[16'h0F0A] <= 180;
        weight_mem[16'h0F0B] <= 176;
        weight_mem[16'h0F0C] <= 168;
        weight_mem[16'h0F0D] <= 162;
        weight_mem[16'h0F0E] <= 155;
        weight_mem[16'h0F0F] <= 146;
        weight_mem[16'h0F10] <= 146;
        weight_mem[16'h0F11] <= 150;
        weight_mem[16'h0F12] <= 156;
        weight_mem[16'h0F13] <= 168;
        weight_mem[16'h0F14] <= 192;
        weight_mem[16'h0F15] <= 215;
        weight_mem[16'h0F16] <= 191;
        weight_mem[16'h0F17] <= 164;
        weight_mem[16'h0F18] <= 151;
        weight_mem[16'h0F19] <= 149;
        weight_mem[16'h0F1A] <= 172;
        weight_mem[16'h0F1B] <= 188;
        weight_mem[16'h0F1C] <= 188;
        weight_mem[16'h0F1D] <= 184;
        weight_mem[16'h0F1E] <= 180;
        weight_mem[16'h0F1F] <= 180;
        weight_mem[16'h0F20] <= 180;
        weight_mem[16'h0F21] <= 180;
        weight_mem[16'h0F22] <= 180;
        weight_mem[16'h0F23] <= 179;
        weight_mem[16'h0F24] <= 175;
        weight_mem[16'h0F25] <= 167;
        weight_mem[16'h0F26] <= 163;
        weight_mem[16'h0F27] <= 154;
        weight_mem[16'h0F28] <= 154;
        weight_mem[16'h0F29] <= 159;
        weight_mem[16'h0F2A] <= 173;
        weight_mem[16'h0F2B] <= 175;
        weight_mem[16'h0F2C] <= 188;
        weight_mem[16'h0F2D] <= 198;
        weight_mem[16'h0F2E] <= 170;
        weight_mem[16'h0F2F] <= 158;
        weight_mem[16'h0F30] <= 152;
        weight_mem[16'h0F31] <= 156;
        weight_mem[16'h0F32] <= 170;
        weight_mem[16'h0F33] <= 183;
        weight_mem[16'h0F34] <= 188;
        weight_mem[16'h0F35] <= 186;
        weight_mem[16'h0F36] <= 181;
        weight_mem[16'h0F37] <= 180;
        weight_mem[16'h0F38] <= 180;
        weight_mem[16'h0F39] <= 180;
        weight_mem[16'h0F3A] <= 180;
        weight_mem[16'h0F3B] <= 178;
        weight_mem[16'h0F3C] <= 174;
        weight_mem[16'h0F3D] <= 169;
        weight_mem[16'h0F3E] <= 167;
        weight_mem[16'h0F3F] <= 168;
        weight_mem[16'h0F40] <= 170;
        weight_mem[16'h0F41] <= 175;
        weight_mem[16'h0F42] <= 183;
        weight_mem[16'h0F43] <= 172;
        weight_mem[16'h0F44] <= 154;
        weight_mem[16'h0F45] <= 154;
        weight_mem[16'h0F46] <= 147;
        weight_mem[16'h0F47] <= 154;
        weight_mem[16'h0F48] <= 170;
        weight_mem[16'h0F49] <= 169;
        weight_mem[16'h0F4A] <= 174;
        weight_mem[16'h0F4B] <= 179;
        weight_mem[16'h0F4C] <= 182;
        weight_mem[16'h0F4D] <= 183;
        weight_mem[16'h0F4E] <= 181;
        weight_mem[16'h0F4F] <= 180;
        weight_mem[16'h0F50] <= 180;
        weight_mem[16'h0F51] <= 180;
        weight_mem[16'h0F52] <= 179;
        weight_mem[16'h0F53] <= 174;
        weight_mem[16'h0F54] <= 167;
        weight_mem[16'h0F55] <= 162;
        weight_mem[16'h0F56] <= 165;
        weight_mem[16'h0F57] <= 171;
        weight_mem[16'h0F58] <= 157;
        weight_mem[16'h0F59] <= 163;
        weight_mem[16'h0F5A] <= 167;
        weight_mem[16'h0F5B] <= 156;
        weight_mem[16'h0F5C] <= 154;
        weight_mem[16'h0F5D] <= 158;
        weight_mem[16'h0F5E] <= 166;
        weight_mem[16'h0F5F] <= 172;
        weight_mem[16'h0F60] <= 175;
        weight_mem[16'h0F61] <= 176;
        weight_mem[16'h0F62] <= 176;
        weight_mem[16'h0F63] <= 177;
        weight_mem[16'h0F64] <= 179;
        weight_mem[16'h0F65] <= 180;
        weight_mem[16'h0F66] <= 180;
        weight_mem[16'h0F67] <= 180;
        weight_mem[16'h0F68] <= 180;
        weight_mem[16'h0F69] <= 180;
        weight_mem[16'h0F6A] <= 178;
        weight_mem[16'h0F6B] <= 174;
        weight_mem[16'h0F6C] <= 171;
        weight_mem[16'h0F6D] <= 169;
        weight_mem[16'h0F6E] <= 172;
        weight_mem[16'h0F6F] <= 184;
        weight_mem[16'h0F70] <= 185;
        weight_mem[16'h0F71] <= 181;
        weight_mem[16'h0F72] <= 190;
        weight_mem[16'h0F73] <= 190;
        weight_mem[16'h0F74] <= 189;
        weight_mem[16'h0F75] <= 187;
        weight_mem[16'h0F76] <= 190;
        weight_mem[16'h0F77] <= 186;
        weight_mem[16'h0F78] <= 179;
        weight_mem[16'h0F79] <= 178;
        weight_mem[16'h0F7A] <= 180;
        weight_mem[16'h0F7B] <= 178;
        weight_mem[16'h0F7C] <= 179;
        weight_mem[16'h0F7D] <= 180;
        weight_mem[16'h0F7E] <= 180;
        weight_mem[16'h0F7F] <= 180;
        weight_mem[16'h0F80] <= 180;
        weight_mem[16'h0F81] <= 180;
        weight_mem[16'h0F82] <= 179;
        weight_mem[16'h0F83] <= 179;
        weight_mem[16'h0F84] <= 179;
        weight_mem[16'h0F85] <= 178;
        weight_mem[16'h0F86] <= 180;
        weight_mem[16'h0F87] <= 186;
        weight_mem[16'h0F88] <= 193;
        weight_mem[16'h0F89] <= 195;
        weight_mem[16'h0F8A] <= 195;
        weight_mem[16'h0F8B] <= 188;
        weight_mem[16'h0F8C] <= 187;
        weight_mem[16'h0F8D] <= 188;
        weight_mem[16'h0F8E] <= 185;
        weight_mem[16'h0F8F] <= 181;
        weight_mem[16'h0F90] <= 179;
        weight_mem[16'h0F91] <= 178;
        weight_mem[16'h0F92] <= 179;
        weight_mem[16'h0F93] <= 179;
        weight_mem[16'h0F94] <= 179;
        weight_mem[16'h0F95] <= 180;
        weight_mem[16'h0F96] <= 180;
        weight_mem[16'h0F97] <= 180;
        weight_mem[16'h0F98] <= 180;
        weight_mem[16'h0F99] <= 180;
        weight_mem[16'h0F9A] <= 180;
        weight_mem[16'h0F9B] <= 180;
        weight_mem[16'h0F9C] <= 180;
        weight_mem[16'h0F9D] <= 180;
        weight_mem[16'h0F9E] <= 180;
        weight_mem[16'h0F9F] <= 180;
        weight_mem[16'h0FA0] <= 182;
        weight_mem[16'h0FA1] <= 183;
        weight_mem[16'h0FA2] <= 182;
        weight_mem[16'h0FA3] <= 181;
        weight_mem[16'h0FA4] <= 182;
        weight_mem[16'h0FA5] <= 182;
        weight_mem[16'h0FA6] <= 180;
        weight_mem[16'h0FA7] <= 180;
        weight_mem[16'h0FA8] <= 180;
        weight_mem[16'h0FA9] <= 179;
        weight_mem[16'h0FAA] <= 179;
        weight_mem[16'h0FAB] <= 180;
        weight_mem[16'h0FAC] <= 180;
        weight_mem[16'h0FAD] <= 180;
        weight_mem[16'h0FAE] <= 180;
        weight_mem[16'h0FAF] <= 180;

        // layer 1 neuron 8
        weight_mem[16'h1000] <= 11;
        weight_mem[16'h1001] <= 4;
        weight_mem[16'h1002] <= 12;
        weight_mem[16'h1003] <= 6;
        weight_mem[16'h1004] <= 11;
        weight_mem[16'h1005] <= 6;
        weight_mem[16'h1006] <= 11;
        weight_mem[16'h1007] <= 11;
        weight_mem[16'h1008] <= 7;
        weight_mem[16'h1009] <= 0;
        weight_mem[16'h100A] <= 5;
        weight_mem[16'h100B] <= 12;
        weight_mem[16'h100C] <= 11;
        weight_mem[16'h100D] <= 4;
        weight_mem[16'h100E] <= 7;
        weight_mem[16'h100F] <= 0;
        weight_mem[16'h1010] <= 10;
        weight_mem[16'h1011] <= 8;
        weight_mem[16'h1012] <= 5;
        weight_mem[16'h1013] <= 13;
        weight_mem[16'h1014] <= 13;
        weight_mem[16'h1015] <= 10;
        weight_mem[16'h1016] <= 1;
        weight_mem[16'h1017] <= 255;
        weight_mem[16'h1018] <= 254;
        weight_mem[16'h1019] <= 253;
        weight_mem[16'h101A] <= 10;
        weight_mem[16'h101B] <= 11;
        weight_mem[16'h101C] <= 5;
        weight_mem[16'h101D] <= 12;
        weight_mem[16'h101E] <= 12;
        weight_mem[16'h101F] <= 3;
        weight_mem[16'h1020] <= 252;
        weight_mem[16'h1021] <= 2;
        weight_mem[16'h1022] <= 10;
        weight_mem[16'h1023] <= 8;
        weight_mem[16'h1024] <= 9;
        weight_mem[16'h1025] <= 254;
        weight_mem[16'h1026] <= 6;
        weight_mem[16'h1027] <= 0;
        weight_mem[16'h1028] <= 4;
        weight_mem[16'h1029] <= 0;
        weight_mem[16'h102A] <= 12;
        weight_mem[16'h102B] <= 6;
        weight_mem[16'h102C] <= 6;
        weight_mem[16'h102D] <= 255;
        weight_mem[16'h102E] <= 7;
        weight_mem[16'h102F] <= 11;
        weight_mem[16'h1030] <= 9;
        weight_mem[16'h1031] <= 254;
        weight_mem[16'h1032] <= 7;
        weight_mem[16'h1033] <= 5;
        weight_mem[16'h1034] <= 12;
        weight_mem[16'h1035] <= 11;
        weight_mem[16'h1036] <= 0;
        weight_mem[16'h1037] <= 3;
        weight_mem[16'h1038] <= 0;
        weight_mem[16'h1039] <= 252;
        weight_mem[16'h103A] <= 4;
        weight_mem[16'h103B] <= 4;
        weight_mem[16'h103C] <= 252;
        weight_mem[16'h103D] <= 12;
        weight_mem[16'h103E] <= 1;
        weight_mem[16'h103F] <= 0;
        weight_mem[16'h1040] <= 10;
        weight_mem[16'h1041] <= 254;
        weight_mem[16'h1042] <= 0;
        weight_mem[16'h1043] <= 255;
        weight_mem[16'h1044] <= 7;
        weight_mem[16'h1045] <= 4;
        weight_mem[16'h1046] <= 9;
        weight_mem[16'h1047] <= 3;
        weight_mem[16'h1048] <= 254;
        weight_mem[16'h1049] <= 4;
        weight_mem[16'h104A] <= 0;
        weight_mem[16'h104B] <= 2;
        weight_mem[16'h104C] <= 4;
        weight_mem[16'h104D] <= 3;
        weight_mem[16'h104E] <= 6;
        weight_mem[16'h104F] <= 253;
        weight_mem[16'h1050] <= 254;
        weight_mem[16'h1051] <= 248;
        weight_mem[16'h1052] <= 248;
        weight_mem[16'h1053] <= 244;
        weight_mem[16'h1054] <= 255;
        weight_mem[16'h1055] <= 253;
        weight_mem[16'h1056] <= 246;
        weight_mem[16'h1057] <= 4;
        weight_mem[16'h1058] <= 248;
        weight_mem[16'h1059] <= 243;
        weight_mem[16'h105A] <= 255;
        weight_mem[16'h105B] <= 2;
        weight_mem[16'h105C] <= 251;
        weight_mem[16'h105D] <= 250;
        weight_mem[16'h105E] <= 252;
        weight_mem[16'h105F] <= 2;
        weight_mem[16'h1060] <= 6;
        weight_mem[16'h1061] <= 9;
        weight_mem[16'h1062] <= 9;
        weight_mem[16'h1063] <= 13;
        weight_mem[16'h1064] <= 13;
        weight_mem[16'h1065] <= 13;
        weight_mem[16'h1066] <= 5;
        weight_mem[16'h1067] <= 6;
        weight_mem[16'h1068] <= 4;
        weight_mem[16'h1069] <= 0;
        weight_mem[16'h106A] <= 236;
        weight_mem[16'h106B] <= 231;
        weight_mem[16'h106C] <= 231;
        weight_mem[16'h106D] <= 222;
        weight_mem[16'h106E] <= 249;
        weight_mem[16'h106F] <= 5;
        weight_mem[16'h1070] <= 2;
        weight_mem[16'h1071] <= 0;
        weight_mem[16'h1072] <= 250;
        weight_mem[16'h1073] <= 244;
        weight_mem[16'h1074] <= 231;
        weight_mem[16'h1075] <= 246;
        weight_mem[16'h1076] <= 248;
        weight_mem[16'h1077] <= 255;
        weight_mem[16'h1078] <= 10;
        weight_mem[16'h1079] <= 1;
        weight_mem[16'h107A] <= 7;
        weight_mem[16'h107B] <= 15;
        weight_mem[16'h107C] <= 14;
        weight_mem[16'h107D] <= 4;
        weight_mem[16'h107E] <= 2;
        weight_mem[16'h107F] <= 242;
        weight_mem[16'h1080] <= 230;
        weight_mem[16'h1081] <= 219;
        weight_mem[16'h1082] <= 195;
        weight_mem[16'h1083] <= 192;
        weight_mem[16'h1084] <= 225;
        weight_mem[16'h1085] <= 1;
        weight_mem[16'h1086] <= 7;
        weight_mem[16'h1087] <= 0;
        weight_mem[16'h1088] <= 0;
        weight_mem[16'h1089] <= 251;
        weight_mem[16'h108A] <= 251;
        weight_mem[16'h108B] <= 252;
        weight_mem[16'h108C] <= 233;
        weight_mem[16'h108D] <= 230;
        weight_mem[16'h108E] <= 247;
        weight_mem[16'h108F] <= 6;
        weight_mem[16'h1090] <= 254;
        weight_mem[16'h1091] <= 3;
        weight_mem[16'h1092] <= 7;
        weight_mem[16'h1093] <= 11;
        weight_mem[16'h1094] <= 4;
        weight_mem[16'h1095] <= 246;
        weight_mem[16'h1096] <= 244;
        weight_mem[16'h1097] <= 230;
        weight_mem[16'h1098] <= 213;
        weight_mem[16'h1099] <= 213;
        weight_mem[16'h109A] <= 227;
        weight_mem[16'h109B] <= 9;
        weight_mem[16'h109C] <= 35;
        weight_mem[16'h109D] <= 49;
        weight_mem[16'h109E] <= 44;
        weight_mem[16'h109F] <= 25;
        weight_mem[16'h10A0] <= 24;
        weight_mem[16'h10A1] <= 32;
        weight_mem[16'h10A2] <= 27;
        weight_mem[16'h10A3] <= 13;
        weight_mem[16'h10A4] <= 0;
        weight_mem[16'h10A5] <= 241;
        weight_mem[16'h10A6] <= 253;
        weight_mem[16'h10A7] <= 254;
        weight_mem[16'h10A8] <= 255;
        weight_mem[16'h10A9] <= 8;
        weight_mem[16'h10AA] <= 9;
        weight_mem[16'h10AB] <= 9;
        weight_mem[16'h10AC] <= 7;
        weight_mem[16'h10AD] <= 247;
        weight_mem[16'h10AE] <= 251;
        weight_mem[16'h10AF] <= 246;
        weight_mem[16'h10B0] <= 233;
        weight_mem[16'h10B1] <= 1;
        weight_mem[16'h10B2] <= 28;
        weight_mem[16'h10B3] <= 23;
        weight_mem[16'h10B4] <= 12;
        weight_mem[16'h10B5] <= 31;
        weight_mem[16'h10B6] <= 47;
        weight_mem[16'h10B7] <= 39;
        weight_mem[16'h10B8] <= 31;
        weight_mem[16'h10B9] <= 24;
        weight_mem[16'h10BA] <= 45;
        weight_mem[16'h10BB] <= 39;
        weight_mem[16'h10BC] <= 20;
        weight_mem[16'h10BD] <= 1;
        weight_mem[16'h10BE] <= 247;
        weight_mem[16'h10BF] <= 7;
        weight_mem[16'h10C0] <= 1;
        weight_mem[16'h10C1] <= 5;
        weight_mem[16'h10C2] <= 10;
        weight_mem[16'h10C3] <= 10;
        weight_mem[16'h10C4] <= 20;
        weight_mem[16'h10C5] <= 23;
        weight_mem[16'h10C6] <= 6;
        weight_mem[16'h10C7] <= 4;
        weight_mem[16'h10C8] <= 19;
        weight_mem[16'h10C9] <= 33;
        weight_mem[16'h10CA] <= 23;
        weight_mem[16'h10CB] <= 234;
        weight_mem[16'h10CC] <= 218;
        weight_mem[16'h10CD] <= 237;
        weight_mem[16'h10CE] <= 10;
        weight_mem[16'h10CF] <= 9;
        weight_mem[16'h10D0] <= 3;
        weight_mem[16'h10D1] <= 3;
        weight_mem[16'h10D2] <= 41;
        weight_mem[16'h10D3] <= 54;
        weight_mem[16'h10D4] <= 41;
        weight_mem[16'h10D5] <= 5;
        weight_mem[16'h10D6] <= 252;
        weight_mem[16'h10D7] <= 11;
        weight_mem[16'h10D8] <= 0;
        weight_mem[16'h10D9] <= 1;
        weight_mem[16'h10DA] <= 10;
        weight_mem[16'h10DB] <= 2;
        weight_mem[16'h10DC] <= 29;
        weight_mem[16'h10DD] <= 32;
        weight_mem[16'h10DE] <= 25;
        weight_mem[16'h10DF] <= 14;
        weight_mem[16'h10E0] <= 24;
        weight_mem[16'h10E1] <= 29;
        weight_mem[16'h10E2] <= 237;
        weight_mem[16'h10E3] <= 185;
        weight_mem[16'h10E4] <= 177;
        weight_mem[16'h10E5] <= 222;
        weight_mem[16'h10E6] <= 3;
        weight_mem[16'h10E7] <= 8;
        weight_mem[16'h10E8] <= 14;
        weight_mem[16'h10E9] <= 35;
        weight_mem[16'h10EA] <= 43;
        weight_mem[16'h10EB] <= 53;
        weight_mem[16'h10EC] <= 38;
        weight_mem[16'h10ED] <= 4;
        weight_mem[16'h10EE] <= 255;
        weight_mem[16'h10EF] <= 7;
        weight_mem[16'h10F0] <= 13;
        weight_mem[16'h10F1] <= 4;
        weight_mem[16'h10F2] <= 6;
        weight_mem[16'h10F3] <= 8;
        weight_mem[16'h10F4] <= 26;
        weight_mem[16'h10F5] <= 19;
        weight_mem[16'h10F6] <= 25;
        weight_mem[16'h10F7] <= 12;
        weight_mem[16'h10F8] <= 9;
        weight_mem[16'h10F9] <= 250;
        weight_mem[16'h10FA] <= 175;
        weight_mem[16'h10FB] <= 128;
        weight_mem[16'h10FC] <= 145;
        weight_mem[16'h10FD] <= 218;
        weight_mem[16'h10FE] <= 0;
        weight_mem[16'h10FF] <= 24;
        weight_mem[16'h1100] <= 35;
        weight_mem[16'h1101] <= 42;
        weight_mem[16'h1102] <= 33;
        weight_mem[16'h1103] <= 29;
        weight_mem[16'h1104] <= 20;
        weight_mem[16'h1105] <= 1;
        weight_mem[16'h1106] <= 251;
        weight_mem[16'h1107] <= 1;
        weight_mem[16'h1108] <= 9;
        weight_mem[16'h1109] <= 12;
        weight_mem[16'h110A] <= 250;
        weight_mem[16'h110B] <= 7;
        weight_mem[16'h110C] <= 12;
        weight_mem[16'h110D] <= 255;
        weight_mem[16'h110E] <= 10;
        weight_mem[16'h110F] <= 0;
        weight_mem[16'h1110] <= 0;
        weight_mem[16'h1111] <= 227;
        weight_mem[16'h1112] <= 185;
        weight_mem[16'h1113] <= 168;
        weight_mem[16'h1114] <= 201;
        weight_mem[16'h1115] <= 248;
        weight_mem[16'h1116] <= 22;
        weight_mem[16'h1117] <= 31;
        weight_mem[16'h1118] <= 10;
        weight_mem[16'h1119] <= 8;
        weight_mem[16'h111A] <= 12;
        weight_mem[16'h111B] <= 5;
        weight_mem[16'h111C] <= 243;
        weight_mem[16'h111D] <= 241;
        weight_mem[16'h111E] <= 0;
        weight_mem[16'h111F] <= 5;
        weight_mem[16'h1120] <= 13;
        weight_mem[16'h1121] <= 10;
        weight_mem[16'h1122] <= 251;
        weight_mem[16'h1123] <= 3;
        weight_mem[16'h1124] <= 3;
        weight_mem[16'h1125] <= 246;
        weight_mem[16'h1126] <= 229;
        weight_mem[16'h1127] <= 244;
        weight_mem[16'h1128] <= 251;
        weight_mem[16'h1129] <= 5;
        weight_mem[16'h112A] <= 245;
        weight_mem[16'h112B] <= 232;
        weight_mem[16'h112C] <= 242;
        weight_mem[16'h112D] <= 7;
        weight_mem[16'h112E] <= 19;
        weight_mem[16'h112F] <= 3;
        weight_mem[16'h1130] <= 5;
        weight_mem[16'h1131] <= 241;
        weight_mem[16'h1132] <= 234;
        weight_mem[16'h1133] <= 227;
        weight_mem[16'h1134] <= 236;
        weight_mem[16'h1135] <= 254;
        weight_mem[16'h1136] <= 10;
        weight_mem[16'h1137] <= 0;
        weight_mem[16'h1138] <= 9;
        weight_mem[16'h1139] <= 3;
        weight_mem[16'h113A] <= 255;
        weight_mem[16'h113B] <= 250;
        weight_mem[16'h113C] <= 3;
        weight_mem[16'h113D] <= 246;
        weight_mem[16'h113E] <= 231;
        weight_mem[16'h113F] <= 232;
        weight_mem[16'h1140] <= 237;
        weight_mem[16'h1141] <= 7;
        weight_mem[16'h1142] <= 11;
        weight_mem[16'h1143] <= 8;
        weight_mem[16'h1144] <= 21;
        weight_mem[16'h1145] <= 26;
        weight_mem[16'h1146] <= 24;
        weight_mem[16'h1147] <= 8;
        weight_mem[16'h1148] <= 244;
        weight_mem[16'h1149] <= 231;
        weight_mem[16'h114A] <= 229;
        weight_mem[16'h114B] <= 222;
        weight_mem[16'h114C] <= 243;
        weight_mem[16'h114D] <= 4;
        weight_mem[16'h114E] <= 7;
        weight_mem[16'h114F] <= 0;
        weight_mem[16'h1150] <= 254;
        weight_mem[16'h1151] <= 0;
        weight_mem[16'h1152] <= 12;
        weight_mem[16'h1153] <= 2;
        weight_mem[16'h1154] <= 4;
        weight_mem[16'h1155] <= 253;
        weight_mem[16'h1156] <= 8;
        weight_mem[16'h1157] <= 253;
        weight_mem[16'h1158] <= 247;
        weight_mem[16'h1159] <= 253;
        weight_mem[16'h115A] <= 15;
        weight_mem[16'h115B] <= 15;
        weight_mem[16'h115C] <= 26;
        weight_mem[16'h115D] <= 20;
        weight_mem[16'h115E] <= 1;
        weight_mem[16'h115F] <= 234;
        weight_mem[16'h1160] <= 216;
        weight_mem[16'h1161] <= 215;
        weight_mem[16'h1162] <= 225;
        weight_mem[16'h1163] <= 247;
        weight_mem[16'h1164] <= 1;
        weight_mem[16'h1165] <= 253;
        weight_mem[16'h1166] <= 0;
        weight_mem[16'h1167] <= 0;
        weight_mem[16'h1168] <= 0;
        weight_mem[16'h1169] <= 254;
        weight_mem[16'h116A] <= 2;
        weight_mem[16'h116B] <= 7;
        weight_mem[16'h116C] <= 16;
        weight_mem[16'h116D] <= 19;
        weight_mem[16'h116E] <= 23;
        weight_mem[16'h116F] <= 13;
        weight_mem[16'h1170] <= 1;
        weight_mem[16'h1171] <= 14;
        weight_mem[16'h1172] <= 248;
        weight_mem[16'h1173] <= 252;
        weight_mem[16'h1174] <= 0;
        weight_mem[16'h1175] <= 249;
        weight_mem[16'h1176] <= 238;
        weight_mem[16'h1177] <= 240;
        weight_mem[16'h1178] <= 237;
        weight_mem[16'h1179] <= 244;
        weight_mem[16'h117A] <= 242;
        weight_mem[16'h117B] <= 252;
        weight_mem[16'h117C] <= 252;
        weight_mem[16'h117D] <= 2;
        weight_mem[16'h117E] <= 9;
        weight_mem[16'h117F] <= 0;
        weight_mem[16'h1180] <= 11;
        weight_mem[16'h1181] <= 5;
        weight_mem[16'h1182] <= 10;
        weight_mem[16'h1183] <= 3;
        weight_mem[16'h1184] <= 7;
        weight_mem[16'h1185] <= 17;
        weight_mem[16'h1186] <= 14;
        weight_mem[16'h1187] <= 16;
        weight_mem[16'h1188] <= 8;
        weight_mem[16'h1189] <= 11;
        weight_mem[16'h118A] <= 5;
        weight_mem[16'h118B] <= 1;
        weight_mem[16'h118C] <= 252;
        weight_mem[16'h118D] <= 253;
        weight_mem[16'h118E] <= 2;
        weight_mem[16'h118F] <= 250;
        weight_mem[16'h1190] <= 248;
        weight_mem[16'h1191] <= 246;
        weight_mem[16'h1192] <= 249;
        weight_mem[16'h1193] <= 9;
        weight_mem[16'h1194] <= 7;
        weight_mem[16'h1195] <= 7;
        weight_mem[16'h1196] <= 13;
        weight_mem[16'h1197] <= 11;
        weight_mem[16'h1198] <= 10;
        weight_mem[16'h1199] <= 254;
        weight_mem[16'h119A] <= 255;
        weight_mem[16'h119B] <= 5;
        weight_mem[16'h119C] <= 4;
        weight_mem[16'h119D] <= 0;
        weight_mem[16'h119E] <= 5;
        weight_mem[16'h119F] <= 13;
        weight_mem[16'h11A0] <= 2;
        weight_mem[16'h11A1] <= 0;
        weight_mem[16'h11A2] <= 2;
        weight_mem[16'h11A3] <= 12;
        weight_mem[16'h11A4] <= 11;
        weight_mem[16'h11A5] <= 10;
        weight_mem[16'h11A6] <= 8;
        weight_mem[16'h11A7] <= 15;
        weight_mem[16'h11A8] <= 5;
        weight_mem[16'h11A9] <= 0;
        weight_mem[16'h11AA] <= 253;
        weight_mem[16'h11AB] <= 6;
        weight_mem[16'h11AC] <= 7;
        weight_mem[16'h11AD] <= 11;
        weight_mem[16'h11AE] <= 13;
        weight_mem[16'h11AF] <= 10;

        // layer 1 neuron 9
        weight_mem[16'h1200] <= 251;
        weight_mem[16'h1201] <= 13;
        weight_mem[16'h1202] <= 6;
        weight_mem[16'h1203] <= 250;
        weight_mem[16'h1204] <= 15;
        weight_mem[16'h1205] <= 8;
        weight_mem[16'h1206] <= 16;
        weight_mem[16'h1207] <= 250;
        weight_mem[16'h1208] <= 13;
        weight_mem[16'h1209] <= 5;
        weight_mem[16'h120A] <= 0;
        weight_mem[16'h120B] <= 13;
        weight_mem[16'h120C] <= 15;
        weight_mem[16'h120D] <= 250;
        weight_mem[16'h120E] <= 254;
        weight_mem[16'h120F] <= 15;
        weight_mem[16'h1210] <= 13;
        weight_mem[16'h1211] <= 7;
        weight_mem[16'h1212] <= 254;
        weight_mem[16'h1213] <= 15;
        weight_mem[16'h1214] <= 4;
        weight_mem[16'h1215] <= 252;
        weight_mem[16'h1216] <= 16;
        weight_mem[16'h1217] <= 17;
        weight_mem[16'h1218] <= 8;
        weight_mem[16'h1219] <= 19;
        weight_mem[16'h121A] <= 7;
        weight_mem[16'h121B] <= 12;
        weight_mem[16'h121C] <= 10;
        weight_mem[16'h121D] <= 5;
        weight_mem[16'h121E] <= 2;
        weight_mem[16'h121F] <= 11;
        weight_mem[16'h1220] <= 249;
        weight_mem[16'h1221] <= 10;
        weight_mem[16'h1222] <= 246;
        weight_mem[16'h1223] <= 6;
        weight_mem[16'h1224] <= 246;
        weight_mem[16'h1225] <= 5;
        weight_mem[16'h1226] <= 254;
        weight_mem[16'h1227] <= 15;
        weight_mem[16'h1228] <= 17;
        weight_mem[16'h1229] <= 13;
        weight_mem[16'h122A] <= 9;
        weight_mem[16'h122B] <= 11;
        weight_mem[16'h122C] <= 10;
        weight_mem[16'h122D] <= 254;
        weight_mem[16'h122E] <= 4;
        weight_mem[16'h122F] <= 0;
        weight_mem[16'h1230] <= 253;
        weight_mem[16'h1231] <= 14;
        weight_mem[16'h1232] <= 4;
        weight_mem[16'h1233] <= 16;
        weight_mem[16'h1234] <= 2;
        weight_mem[16'h1235] <= 12;
        weight_mem[16'h1236] <= 244;
        weight_mem[16'h1237] <= 238;
        weight_mem[16'h1238] <= 223;
        weight_mem[16'h1239] <= 207;
        weight_mem[16'h123A] <= 203;
        weight_mem[16'h123B] <= 212;
        weight_mem[16'h123C] <= 227;
        weight_mem[16'h123D] <= 227;
        weight_mem[16'h123E] <= 1;
        weight_mem[16'h123F] <= 247;
        weight_mem[16'h1240] <= 12;
        weight_mem[16'h1241] <= 20;
        weight_mem[16'h1242] <= 27;
        weight_mem[16'h1243] <= 21;
        weight_mem[16'h1244] <= 22;
        weight_mem[16'h1245] <= 15;
        weight_mem[16'h1246] <= 8;
        weight_mem[16'h1247] <= 252;
        weight_mem[16'h1248] <= 1;
        weight_mem[16'h1249] <= 3;
        weight_mem[16'h124A] <= 10;
        weight_mem[16'h124B] <= 248;
        weight_mem[16'h124C] <= 247;
        weight_mem[16'h124D] <= 245;
        weight_mem[16'h124E] <= 224;
        weight_mem[16'h124F] <= 206;
        weight_mem[16'h1250] <= 193;
        weight_mem[16'h1251] <= 197;
        weight_mem[16'h1252] <= 203;
        weight_mem[16'h1253] <= 201;
        weight_mem[16'h1254] <= 209;
        weight_mem[16'h1255] <= 207;
        weight_mem[16'h1256] <= 199;
        weight_mem[16'h1257] <= 228;
        weight_mem[16'h1258] <= 5;
        weight_mem[16'h1259] <= 5;
        weight_mem[16'h125A] <= 34;
        weight_mem[16'h125B] <= 42;
        weight_mem[16'h125C] <= 39;
        weight_mem[16'h125D] <= 13;
        weight_mem[16'h125E] <= 14;
        weight_mem[16'h125F] <= 10;
        weight_mem[16'h1260] <= 7;
        weight_mem[16'h1261] <= 17;
        weight_mem[16'h1262] <= 8;
        weight_mem[16'h1263] <= 244;
        weight_mem[16'h1264] <= 252;
        weight_mem[16'h1265] <= 227;
        weight_mem[16'h1266] <= 227;
        weight_mem[16'h1267] <= 213;
        weight_mem[16'h1268] <= 216;
        weight_mem[16'h1269] <= 215;
        weight_mem[16'h126A] <= 206;
        weight_mem[16'h126B] <= 174;
        weight_mem[16'h126C] <= 175;
        weight_mem[16'h126D] <= 186;
        weight_mem[16'h126E] <= 202;
        weight_mem[16'h126F] <= 211;
        weight_mem[16'h1270] <= 229;
        weight_mem[16'h1271] <= 248;
        weight_mem[16'h1272] <= 2;
        weight_mem[16'h1273] <= 14;
        weight_mem[16'h1274] <= 48;
        weight_mem[16'h1275] <= 31;
        weight_mem[16'h1276] <= 0;
        weight_mem[16'h1277] <= 11;
        weight_mem[16'h1278] <= 250;
        weight_mem[16'h1279] <= 16;
        weight_mem[16'h127A] <= 7;
        weight_mem[16'h127B] <= 252;
        weight_mem[16'h127C] <= 251;
        weight_mem[16'h127D] <= 249;
        weight_mem[16'h127E] <= 252;
        weight_mem[16'h127F] <= 253;
        weight_mem[16'h1280] <= 248;
        weight_mem[16'h1281] <= 219;
        weight_mem[16'h1282] <= 224;
        weight_mem[16'h1283] <= 221;
        weight_mem[16'h1284] <= 184;
        weight_mem[16'h1285] <= 179;
        weight_mem[16'h1286] <= 192;
        weight_mem[16'h1287] <= 205;
        weight_mem[16'h1288] <= 213;
        weight_mem[16'h1289] <= 223;
        weight_mem[16'h128A] <= 234;
        weight_mem[16'h128B] <= 1;
        weight_mem[16'h128C] <= 43;
        weight_mem[16'h128D] <= 21;
        weight_mem[16'h128E] <= 13;
        weight_mem[16'h128F] <= 5;
        weight_mem[16'h1290] <= 8;
        weight_mem[16'h1291] <= 4;
        weight_mem[16'h1292] <= 9;
        weight_mem[16'h1293] <= 0;
        weight_mem[16'h1294] <= 255;
        weight_mem[16'h1295] <= 18;
        weight_mem[16'h1296] <= 44;
        weight_mem[16'h1297] <= 33;
        weight_mem[16'h1298] <= 51;
        weight_mem[16'h1299] <= 66;
        weight_mem[16'h129A] <= 90;
        weight_mem[16'h129B] <= 85;
        weight_mem[16'h129C] <= 28;
        weight_mem[16'h129D] <= 248;
        weight_mem[16'h129E] <= 203;
        weight_mem[16'h129F] <= 216;
        weight_mem[16'h12A0] <= 218;
        weight_mem[16'h12A1] <= 208;
        weight_mem[16'h12A2] <= 212;
        weight_mem[16'h12A3] <= 225;
        weight_mem[16'h12A4] <= 20;
        weight_mem[16'h12A5] <= 17;
        weight_mem[16'h12A6] <= 15;
        weight_mem[16'h12A7] <= 4;
        weight_mem[16'h12A8] <= 17;
        weight_mem[16'h12A9] <= 250;
        weight_mem[16'h12AA] <= 13;
        weight_mem[16'h12AB] <= 2;
        weight_mem[16'h12AC] <= 28;
        weight_mem[16'h12AD] <= 73;
        weight_mem[16'h12AE] <= 65;
        weight_mem[16'h12AF] <= 74;
        weight_mem[16'h12B0] <= 81;
        weight_mem[16'h12B1] <= 79;
        weight_mem[16'h12B2] <= 102;
        weight_mem[16'h12B3] <= 127;
        weight_mem[16'h12B4] <= 93;
        weight_mem[16'h12B5] <= 57;
        weight_mem[16'h12B6] <= 35;
        weight_mem[16'h12B7] <= 245;
        weight_mem[16'h12B8] <= 227;
        weight_mem[16'h12B9] <= 210;
        weight_mem[16'h12BA] <= 233;
        weight_mem[16'h12BB] <= 252;
        weight_mem[16'h12BC] <= 248;
        weight_mem[16'h12BD] <= 255;
        weight_mem[16'h12BE] <= 9;
        weight_mem[16'h12BF] <= 18;
        weight_mem[16'h12C0] <= 5;
        weight_mem[16'h12C1] <= 8;
        weight_mem[16'h12C2] <= 12;
        weight_mem[16'h12C3] <= 19;
        weight_mem[16'h12C4] <= 55;
        weight_mem[16'h12C5] <= 78;
        weight_mem[16'h12C6] <= 63;
        weight_mem[16'h12C7] <= 36;
        weight_mem[16'h12C8] <= 251;
        weight_mem[16'h12C9] <= 243;
        weight_mem[16'h12CA] <= 27;
        weight_mem[16'h12CB] <= 28;
        weight_mem[16'h12CC] <= 55;
        weight_mem[16'h12CD] <= 75;
        weight_mem[16'h12CE] <= 42;
        weight_mem[16'h12CF] <= 11;
        weight_mem[16'h12D0] <= 8;
        weight_mem[16'h12D1] <= 253;
        weight_mem[16'h12D2] <= 21;
        weight_mem[16'h12D3] <= 27;
        weight_mem[16'h12D4] <= 16;
        weight_mem[16'h12D5] <= 14;
        weight_mem[16'h12D6] <= 253;
        weight_mem[16'h12D7] <= 6;
        weight_mem[16'h12D8] <= 11;
        weight_mem[16'h12D9] <= 5;
        weight_mem[16'h12DA] <= 13;
        weight_mem[16'h12DB] <= 18;
        weight_mem[16'h12DC] <= 32;
        weight_mem[16'h12DD] <= 44;
        weight_mem[16'h12DE] <= 251;
        weight_mem[16'h12DF] <= 234;
        weight_mem[16'h12E0] <= 234;
        weight_mem[16'h12E1] <= 244;
        weight_mem[16'h12E2] <= 236;
        weight_mem[16'h12E3] <= 241;
        weight_mem[16'h12E4] <= 1;
        weight_mem[16'h12E5] <= 7;
        weight_mem[16'h12E6] <= 12;
        weight_mem[16'h12E7] <= 250;
        weight_mem[16'h12E8] <= 19;
        weight_mem[16'h12E9] <= 30;
        weight_mem[16'h12EA] <= 34;
        weight_mem[16'h12EB] <= 37;
        weight_mem[16'h12EC] <= 17;
        weight_mem[16'h12ED] <= 255;
        weight_mem[16'h12EE] <= 243;
        weight_mem[16'h12EF] <= 16;
        weight_mem[16'h12F0] <= 6;
        weight_mem[16'h12F1] <= 250;
        weight_mem[16'h12F2] <= 8;
        weight_mem[16'h12F3] <= 241;
        weight_mem[16'h12F4] <= 237;
        weight_mem[16'h12F5] <= 237;
        weight_mem[16'h12F6] <= 3;
        weight_mem[16'h12F7] <= 14;
        weight_mem[16'h12F8] <= 253;
        weight_mem[16'h12F9] <= 7;
        weight_mem[16'h12FA] <= 6;
        weight_mem[16'h12FB] <= 14;
        weight_mem[16'h12FC] <= 18;
        weight_mem[16'h12FD] <= 2;
        weight_mem[16'h12FE] <= 2;
        weight_mem[16'h12FF] <= 5;
        weight_mem[16'h1300] <= 21;
        weight_mem[16'h1301] <= 44;
        weight_mem[16'h1302] <= 23;
        weight_mem[16'h1303] <= 25;
        weight_mem[16'h1304] <= 6;
        weight_mem[16'h1305] <= 245;
        weight_mem[16'h1306] <= 252;
        weight_mem[16'h1307] <= 250;
        weight_mem[16'h1308] <= 18;
        weight_mem[16'h1309] <= 13;
        weight_mem[16'h130A] <= 1;
        weight_mem[16'h130B] <= 231;
        weight_mem[16'h130C] <= 216;
        weight_mem[16'h130D] <= 243;
        weight_mem[16'h130E] <= 0;
        weight_mem[16'h130F] <= 22;
        weight_mem[16'h1310] <= 28;
        weight_mem[16'h1311] <= 24;
        weight_mem[16'h1312] <= 18;
        weight_mem[16'h1313] <= 3;
        weight_mem[16'h1314] <= 28;
        weight_mem[16'h1315] <= 244;
        weight_mem[16'h1316] <= 229;
        weight_mem[16'h1317] <= 4;
        weight_mem[16'h1318] <= 21;
        weight_mem[16'h1319] <= 22;
        weight_mem[16'h131A] <= 5;
        weight_mem[16'h131B] <= 246;
        weight_mem[16'h131C] <= 232;
        weight_mem[16'h131D] <= 223;
        weight_mem[16'h131E] <= 248;
        weight_mem[16'h131F] <= 6;
        weight_mem[16'h1320] <= 16;
        weight_mem[16'h1321] <= 8;
        weight_mem[16'h1322] <= 244;
        weight_mem[16'h1323] <= 231;
        weight_mem[16'h1324] <= 205;
        weight_mem[16'h1325] <= 229;
        weight_mem[16'h1326] <= 239;
        weight_mem[16'h1327] <= 249;
        weight_mem[16'h1328] <= 235;
        weight_mem[16'h1329] <= 232;
        weight_mem[16'h132A] <= 217;
        weight_mem[16'h132B] <= 228;
        weight_mem[16'h132C] <= 245;
        weight_mem[16'h132D] <= 235;
        weight_mem[16'h132E] <= 234;
        weight_mem[16'h132F] <= 0;
        weight_mem[16'h1330] <= 0;
        weight_mem[16'h1331] <= 254;
        weight_mem[16'h1332] <= 248;
        weight_mem[16'h1333] <= 219;
        weight_mem[16'h1334] <= 232;
        weight_mem[16'h1335] <= 244;
        weight_mem[16'h1336] <= 250;
        weight_mem[16'h1337] <= 12;
        weight_mem[16'h1338] <= 252;
        weight_mem[16'h1339] <= 254;
        weight_mem[16'h133A] <= 250;
        weight_mem[16'h133B] <= 218;
        weight_mem[16'h133C] <= 208;
        weight_mem[16'h133D] <= 231;
        weight_mem[16'h133E] <= 230;
        weight_mem[16'h133F] <= 254;
        weight_mem[16'h1340] <= 238;
        weight_mem[16'h1341] <= 242;
        weight_mem[16'h1342] <= 237;
        weight_mem[16'h1343] <= 227;
        weight_mem[16'h1344] <= 253;
        weight_mem[16'h1345] <= 1;
        weight_mem[16'h1346] <= 13;
        weight_mem[16'h1347] <= 255;
        weight_mem[16'h1348] <= 240;
        weight_mem[16'h1349] <= 240;
        weight_mem[16'h134A] <= 220;
        weight_mem[16'h134B] <= 233;
        weight_mem[16'h134C] <= 231;
        weight_mem[16'h134D] <= 242;
        weight_mem[16'h134E] <= 15;
        weight_mem[16'h134F] <= 3;
        weight_mem[16'h1350] <= 12;
        weight_mem[16'h1351] <= 252;
        weight_mem[16'h1352] <= 11;
        weight_mem[16'h1353] <= 248;
        weight_mem[16'h1354] <= 242;
        weight_mem[16'h1355] <= 226;
        weight_mem[16'h1356] <= 240;
        weight_mem[16'h1357] <= 238;
        weight_mem[16'h1358] <= 241;
        weight_mem[16'h1359] <= 235;
        weight_mem[16'h135A] <= 239;
        weight_mem[16'h135B] <= 235;
        weight_mem[16'h135C] <= 239;
        weight_mem[16'h135D] <= 246;
        weight_mem[16'h135E] <= 248;
        weight_mem[16'h135F] <= 255;
        weight_mem[16'h1360] <= 244;
        weight_mem[16'h1361] <= 248;
        weight_mem[16'h1362] <= 252;
        weight_mem[16'h1363] <= 236;
        weight_mem[16'h1364] <= 248;
        weight_mem[16'h1365] <= 250;
        weight_mem[16'h1366] <= 254;
        weight_mem[16'h1367] <= 8;
        weight_mem[16'h1368] <= 16;
        weight_mem[16'h1369] <= 8;
        weight_mem[16'h136A] <= 11;
        weight_mem[16'h136B] <= 14;
        weight_mem[16'h136C] <= 1;
        weight_mem[16'h136D] <= 247;
        weight_mem[16'h136E] <= 250;
        weight_mem[16'h136F] <= 244;
        weight_mem[16'h1370] <= 249;
        weight_mem[16'h1371] <= 250;
        weight_mem[16'h1372] <= 222;
        weight_mem[16'h1373] <= 232;
        weight_mem[16'h1374] <= 227;
        weight_mem[16'h1375] <= 241;
        weight_mem[16'h1376] <= 253;
        weight_mem[16'h1377] <= 0;
        weight_mem[16'h1378] <= 1;
        weight_mem[16'h1379] <= 7;
        weight_mem[16'h137A] <= 3;
        weight_mem[16'h137B] <= 248;
        weight_mem[16'h137C] <= 7;
        weight_mem[16'h137D] <= 6;
        weight_mem[16'h137E] <= 15;
        weight_mem[16'h137F] <= 18;
        weight_mem[16'h1380] <= 14;
        weight_mem[16'h1381] <= 0;
        weight_mem[16'h1382] <= 252;
        weight_mem[16'h1383] <= 6;
        weight_mem[16'h1384] <= 11;
        weight_mem[16'h1385] <= 12;
        weight_mem[16'h1386] <= 3;
        weight_mem[16'h1387] <= 1;
        weight_mem[16'h1388] <= 5;
        weight_mem[16'h1389] <= 231;
        weight_mem[16'h138A] <= 241;
        weight_mem[16'h138B] <= 241;
        weight_mem[16'h138C] <= 229;
        weight_mem[16'h138D] <= 236;
        weight_mem[16'h138E] <= 250;
        weight_mem[16'h138F] <= 251;
        weight_mem[16'h1390] <= 9;
        weight_mem[16'h1391] <= 4;
        weight_mem[16'h1392] <= 4;
        weight_mem[16'h1393] <= 3;
        weight_mem[16'h1394] <= 5;
        weight_mem[16'h1395] <= 14;
        weight_mem[16'h1396] <= 255;
        weight_mem[16'h1397] <= 255;
        weight_mem[16'h1398] <= 4;
        weight_mem[16'h1399] <= 3;
        weight_mem[16'h139A] <= 252;
        weight_mem[16'h139B] <= 15;
        weight_mem[16'h139C] <= 253;
        weight_mem[16'h139D] <= 254;
        weight_mem[16'h139E] <= 1;
        weight_mem[16'h139F] <= 1;
        weight_mem[16'h13A0] <= 250;
        weight_mem[16'h13A1] <= 2;
        weight_mem[16'h13A2] <= 3;
        weight_mem[16'h13A3] <= 253;
        weight_mem[16'h13A4] <= 251;
        weight_mem[16'h13A5] <= 249;
        weight_mem[16'h13A6] <= 15;
        weight_mem[16'h13A7] <= 12;
        weight_mem[16'h13A8] <= 14;
        weight_mem[16'h13A9] <= 14;
        weight_mem[16'h13AA] <= 7;
        weight_mem[16'h13AB] <= 9;
        weight_mem[16'h13AC] <= 6;
        weight_mem[16'h13AD] <= 16;
        weight_mem[16'h13AE] <= 252;
        weight_mem[16'h13AF] <= 251;

        // layer 1 neuron 10
        weight_mem[16'h1400] <= 0;
        weight_mem[16'h1401] <= 0;
        weight_mem[16'h1402] <= 0;
        weight_mem[16'h1403] <= 0;
        weight_mem[16'h1404] <= 0;
        weight_mem[16'h1405] <= 0;
        weight_mem[16'h1406] <= 0;
        weight_mem[16'h1407] <= 0;
        weight_mem[16'h1408] <= 0;
        weight_mem[16'h1409] <= 0;
        weight_mem[16'h140A] <= 0;
        weight_mem[16'h140B] <= 0;
        weight_mem[16'h140C] <= 0;
        weight_mem[16'h140D] <= 0;
        weight_mem[16'h140E] <= 0;
        weight_mem[16'h140F] <= 0;
        weight_mem[16'h1410] <= 0;
        weight_mem[16'h1411] <= 0;
        weight_mem[16'h1412] <= 0;
        weight_mem[16'h1413] <= 0;
        weight_mem[16'h1414] <= 0;
        weight_mem[16'h1415] <= 0;
        weight_mem[16'h1416] <= 0;
        weight_mem[16'h1417] <= 0;
        weight_mem[16'h1418] <= 0;
        weight_mem[16'h1419] <= 0;
        weight_mem[16'h141A] <= 0;
        weight_mem[16'h141B] <= 0;
        weight_mem[16'h141C] <= 0;
        weight_mem[16'h141D] <= 0;
        weight_mem[16'h141E] <= 0;
        weight_mem[16'h141F] <= 0;
        weight_mem[16'h1420] <= 0;
        weight_mem[16'h1421] <= 0;
        weight_mem[16'h1422] <= 0;
        weight_mem[16'h1423] <= 0;
        weight_mem[16'h1424] <= 0;
        weight_mem[16'h1425] <= 0;
        weight_mem[16'h1426] <= 0;
        weight_mem[16'h1427] <= 0;
        weight_mem[16'h1428] <= 0;
        weight_mem[16'h1429] <= 0;
        weight_mem[16'h142A] <= 0;
        weight_mem[16'h142B] <= 0;
        weight_mem[16'h142C] <= 0;
        weight_mem[16'h142D] <= 0;
        weight_mem[16'h142E] <= 0;
        weight_mem[16'h142F] <= 0;
        weight_mem[16'h1430] <= 0;
        weight_mem[16'h1431] <= 0;
        weight_mem[16'h1432] <= 0;
        weight_mem[16'h1433] <= 0;
        weight_mem[16'h1434] <= 0;
        weight_mem[16'h1435] <= 0;
        weight_mem[16'h1436] <= 0;
        weight_mem[16'h1437] <= 0;
        weight_mem[16'h1438] <= 0;
        weight_mem[16'h1439] <= 0;
        weight_mem[16'h143A] <= 0;
        weight_mem[16'h143B] <= 0;
        weight_mem[16'h143C] <= 0;
        weight_mem[16'h143D] <= 0;
        weight_mem[16'h143E] <= 0;
        weight_mem[16'h143F] <= 0;
        weight_mem[16'h1440] <= 0;
        weight_mem[16'h1441] <= 0;
        weight_mem[16'h1442] <= 0;
        weight_mem[16'h1443] <= 0;
        weight_mem[16'h1444] <= 0;
        weight_mem[16'h1445] <= 0;
        weight_mem[16'h1446] <= 0;
        weight_mem[16'h1447] <= 0;
        weight_mem[16'h1448] <= 0;
        weight_mem[16'h1449] <= 0;
        weight_mem[16'h144A] <= 0;
        weight_mem[16'h144B] <= 0;
        weight_mem[16'h144C] <= 0;
        weight_mem[16'h144D] <= 0;
        weight_mem[16'h144E] <= 0;
        weight_mem[16'h144F] <= 0;
        weight_mem[16'h1450] <= 0;
        weight_mem[16'h1451] <= 0;
        weight_mem[16'h1452] <= 0;
        weight_mem[16'h1453] <= 0;
        weight_mem[16'h1454] <= 0;
        weight_mem[16'h1455] <= 0;
        weight_mem[16'h1456] <= 0;
        weight_mem[16'h1457] <= 0;
        weight_mem[16'h1458] <= 0;
        weight_mem[16'h1459] <= 0;
        weight_mem[16'h145A] <= 0;
        weight_mem[16'h145B] <= 0;
        weight_mem[16'h145C] <= 0;
        weight_mem[16'h145D] <= 0;
        weight_mem[16'h145E] <= 0;
        weight_mem[16'h145F] <= 0;
        weight_mem[16'h1460] <= 0;
        weight_mem[16'h1461] <= 0;
        weight_mem[16'h1462] <= 0;
        weight_mem[16'h1463] <= 0;
        weight_mem[16'h1464] <= 0;
        weight_mem[16'h1465] <= 0;
        weight_mem[16'h1466] <= 0;
        weight_mem[16'h1467] <= 0;
        weight_mem[16'h1468] <= 0;
        weight_mem[16'h1469] <= 0;
        weight_mem[16'h146A] <= 0;
        weight_mem[16'h146B] <= 0;
        weight_mem[16'h146C] <= 255;
        weight_mem[16'h146D] <= 0;
        weight_mem[16'h146E] <= 0;
        weight_mem[16'h146F] <= 0;
        weight_mem[16'h1470] <= 0;
        weight_mem[16'h1471] <= 0;
        weight_mem[16'h1472] <= 0;
        weight_mem[16'h1473] <= 0;
        weight_mem[16'h1474] <= 0;
        weight_mem[16'h1475] <= 0;
        weight_mem[16'h1476] <= 0;
        weight_mem[16'h1477] <= 0;
        weight_mem[16'h1478] <= 0;
        weight_mem[16'h1479] <= 0;
        weight_mem[16'h147A] <= 0;
        weight_mem[16'h147B] <= 0;
        weight_mem[16'h147C] <= 0;
        weight_mem[16'h147D] <= 0;
        weight_mem[16'h147E] <= 0;
        weight_mem[16'h147F] <= 0;
        weight_mem[16'h1480] <= 0;
        weight_mem[16'h1481] <= 0;
        weight_mem[16'h1482] <= 0;
        weight_mem[16'h1483] <= 0;
        weight_mem[16'h1484] <= 0;
        weight_mem[16'h1485] <= 0;
        weight_mem[16'h1486] <= 0;
        weight_mem[16'h1487] <= 0;
        weight_mem[16'h1488] <= 0;
        weight_mem[16'h1489] <= 0;
        weight_mem[16'h148A] <= 0;
        weight_mem[16'h148B] <= 0;
        weight_mem[16'h148C] <= 0;
        weight_mem[16'h148D] <= 0;
        weight_mem[16'h148E] <= 0;
        weight_mem[16'h148F] <= 0;
        weight_mem[16'h1490] <= 0;
        weight_mem[16'h1491] <= 0;
        weight_mem[16'h1492] <= 0;
        weight_mem[16'h1493] <= 0;
        weight_mem[16'h1494] <= 0;
        weight_mem[16'h1495] <= 0;
        weight_mem[16'h1496] <= 0;
        weight_mem[16'h1497] <= 0;
        weight_mem[16'h1498] <= 0;
        weight_mem[16'h1499] <= 0;
        weight_mem[16'h149A] <= 0;
        weight_mem[16'h149B] <= 0;
        weight_mem[16'h149C] <= 0;
        weight_mem[16'h149D] <= 0;
        weight_mem[16'h149E] <= 0;
        weight_mem[16'h149F] <= 0;
        weight_mem[16'h14A0] <= 0;
        weight_mem[16'h14A1] <= 0;
        weight_mem[16'h14A2] <= 0;
        weight_mem[16'h14A3] <= 0;
        weight_mem[16'h14A4] <= 0;
        weight_mem[16'h14A5] <= 0;
        weight_mem[16'h14A6] <= 0;
        weight_mem[16'h14A7] <= 0;
        weight_mem[16'h14A8] <= 0;
        weight_mem[16'h14A9] <= 0;
        weight_mem[16'h14AA] <= 0;
        weight_mem[16'h14AB] <= 0;
        weight_mem[16'h14AC] <= 0;
        weight_mem[16'h14AD] <= 0;
        weight_mem[16'h14AE] <= 0;
        weight_mem[16'h14AF] <= 0;
        weight_mem[16'h14B0] <= 0;
        weight_mem[16'h14B1] <= 0;
        weight_mem[16'h14B2] <= 0;
        weight_mem[16'h14B3] <= 0;
        weight_mem[16'h14B4] <= 0;
        weight_mem[16'h14B5] <= 0;
        weight_mem[16'h14B6] <= 0;
        weight_mem[16'h14B7] <= 0;
        weight_mem[16'h14B8] <= 0;
        weight_mem[16'h14B9] <= 0;
        weight_mem[16'h14BA] <= 0;
        weight_mem[16'h14BB] <= 0;
        weight_mem[16'h14BC] <= 0;
        weight_mem[16'h14BD] <= 0;
        weight_mem[16'h14BE] <= 0;
        weight_mem[16'h14BF] <= 0;
        weight_mem[16'h14C0] <= 0;
        weight_mem[16'h14C1] <= 0;
        weight_mem[16'h14C2] <= 0;
        weight_mem[16'h14C3] <= 0;
        weight_mem[16'h14C4] <= 0;
        weight_mem[16'h14C5] <= 0;
        weight_mem[16'h14C6] <= 0;
        weight_mem[16'h14C7] <= 0;
        weight_mem[16'h14C8] <= 0;
        weight_mem[16'h14C9] <= 0;
        weight_mem[16'h14CA] <= 0;
        weight_mem[16'h14CB] <= 0;
        weight_mem[16'h14CC] <= 0;
        weight_mem[16'h14CD] <= 0;
        weight_mem[16'h14CE] <= 0;
        weight_mem[16'h14CF] <= 0;
        weight_mem[16'h14D0] <= 0;
        weight_mem[16'h14D1] <= 0;
        weight_mem[16'h14D2] <= 253;
        weight_mem[16'h14D3] <= 0;
        weight_mem[16'h14D4] <= 0;
        weight_mem[16'h14D5] <= 0;
        weight_mem[16'h14D6] <= 0;
        weight_mem[16'h14D7] <= 0;
        weight_mem[16'h14D8] <= 0;
        weight_mem[16'h14D9] <= 0;
        weight_mem[16'h14DA] <= 0;
        weight_mem[16'h14DB] <= 0;
        weight_mem[16'h14DC] <= 0;
        weight_mem[16'h14DD] <= 0;
        weight_mem[16'h14DE] <= 0;
        weight_mem[16'h14DF] <= 0;
        weight_mem[16'h14E0] <= 0;
        weight_mem[16'h14E1] <= 0;
        weight_mem[16'h14E2] <= 0;
        weight_mem[16'h14E3] <= 0;
        weight_mem[16'h14E4] <= 0;
        weight_mem[16'h14E5] <= 0;
        weight_mem[16'h14E6] <= 0;
        weight_mem[16'h14E7] <= 0;
        weight_mem[16'h14E8] <= 0;
        weight_mem[16'h14E9] <= 251;
        weight_mem[16'h14EA] <= 251;
        weight_mem[16'h14EB] <= 0;
        weight_mem[16'h14EC] <= 0;
        weight_mem[16'h14ED] <= 0;
        weight_mem[16'h14EE] <= 0;
        weight_mem[16'h14EF] <= 0;
        weight_mem[16'h14F0] <= 0;
        weight_mem[16'h14F1] <= 0;
        weight_mem[16'h14F2] <= 0;
        weight_mem[16'h14F3] <= 0;
        weight_mem[16'h14F4] <= 0;
        weight_mem[16'h14F5] <= 0;
        weight_mem[16'h14F6] <= 0;
        weight_mem[16'h14F7] <= 0;
        weight_mem[16'h14F8] <= 0;
        weight_mem[16'h14F9] <= 0;
        weight_mem[16'h14FA] <= 0;
        weight_mem[16'h14FB] <= 0;
        weight_mem[16'h14FC] <= 0;
        weight_mem[16'h14FD] <= 0;
        weight_mem[16'h14FE] <= 0;
        weight_mem[16'h14FF] <= 0;
        weight_mem[16'h1500] <= 0;
        weight_mem[16'h1501] <= 249;
        weight_mem[16'h1502] <= 253;
        weight_mem[16'h1503] <= 0;
        weight_mem[16'h1504] <= 0;
        weight_mem[16'h1505] <= 0;
        weight_mem[16'h1506] <= 0;
        weight_mem[16'h1507] <= 0;
        weight_mem[16'h1508] <= 0;
        weight_mem[16'h1509] <= 0;
        weight_mem[16'h150A] <= 0;
        weight_mem[16'h150B] <= 0;
        weight_mem[16'h150C] <= 0;
        weight_mem[16'h150D] <= 0;
        weight_mem[16'h150E] <= 254;
        weight_mem[16'h150F] <= 253;
        weight_mem[16'h1510] <= 0;
        weight_mem[16'h1511] <= 0;
        weight_mem[16'h1512] <= 0;
        weight_mem[16'h1513] <= 0;
        weight_mem[16'h1514] <= 0;
        weight_mem[16'h1515] <= 0;
        weight_mem[16'h1516] <= 0;
        weight_mem[16'h1517] <= 0;
        weight_mem[16'h1518] <= 0;
        weight_mem[16'h1519] <= 255;
        weight_mem[16'h151A] <= 255;
        weight_mem[16'h151B] <= 0;
        weight_mem[16'h151C] <= 0;
        weight_mem[16'h151D] <= 0;
        weight_mem[16'h151E] <= 0;
        weight_mem[16'h151F] <= 0;
        weight_mem[16'h1520] <= 0;
        weight_mem[16'h1521] <= 0;
        weight_mem[16'h1522] <= 0;
        weight_mem[16'h1523] <= 0;
        weight_mem[16'h1524] <= 0;
        weight_mem[16'h1525] <= 0;
        weight_mem[16'h1526] <= 0;
        weight_mem[16'h1527] <= 255;
        weight_mem[16'h1528] <= 0;
        weight_mem[16'h1529] <= 0;
        weight_mem[16'h152A] <= 0;
        weight_mem[16'h152B] <= 0;
        weight_mem[16'h152C] <= 0;
        weight_mem[16'h152D] <= 0;
        weight_mem[16'h152E] <= 0;
        weight_mem[16'h152F] <= 254;
        weight_mem[16'h1530] <= 255;
        weight_mem[16'h1531] <= 0;
        weight_mem[16'h1532] <= 0;
        weight_mem[16'h1533] <= 0;
        weight_mem[16'h1534] <= 0;
        weight_mem[16'h1535] <= 0;
        weight_mem[16'h1536] <= 0;
        weight_mem[16'h1537] <= 0;
        weight_mem[16'h1538] <= 0;
        weight_mem[16'h1539] <= 0;
        weight_mem[16'h153A] <= 0;
        weight_mem[16'h153B] <= 0;
        weight_mem[16'h153C] <= 0;
        weight_mem[16'h153D] <= 0;
        weight_mem[16'h153E] <= 0;
        weight_mem[16'h153F] <= 0;
        weight_mem[16'h1540] <= 255;
        weight_mem[16'h1541] <= 255;
        weight_mem[16'h1542] <= 255;
        weight_mem[16'h1543] <= 255;
        weight_mem[16'h1544] <= 0;
        weight_mem[16'h1545] <= 0;
        weight_mem[16'h1546] <= 255;
        weight_mem[16'h1547] <= 0;
        weight_mem[16'h1548] <= 0;
        weight_mem[16'h1549] <= 0;
        weight_mem[16'h154A] <= 0;
        weight_mem[16'h154B] <= 0;
        weight_mem[16'h154C] <= 0;
        weight_mem[16'h154D] <= 0;
        weight_mem[16'h154E] <= 0;
        weight_mem[16'h154F] <= 0;
        weight_mem[16'h1550] <= 0;
        weight_mem[16'h1551] <= 0;
        weight_mem[16'h1552] <= 0;
        weight_mem[16'h1553] <= 0;
        weight_mem[16'h1554] <= 0;
        weight_mem[16'h1555] <= 0;
        weight_mem[16'h1556] <= 0;
        weight_mem[16'h1557] <= 0;
        weight_mem[16'h1558] <= 0;
        weight_mem[16'h1559] <= 0;
        weight_mem[16'h155A] <= 0;
        weight_mem[16'h155B] <= 0;
        weight_mem[16'h155C] <= 0;
        weight_mem[16'h155D] <= 0;
        weight_mem[16'h155E] <= 0;
        weight_mem[16'h155F] <= 0;
        weight_mem[16'h1560] <= 0;
        weight_mem[16'h1561] <= 0;
        weight_mem[16'h1562] <= 0;
        weight_mem[16'h1563] <= 0;
        weight_mem[16'h1564] <= 0;
        weight_mem[16'h1565] <= 0;
        weight_mem[16'h1566] <= 0;
        weight_mem[16'h1567] <= 0;
        weight_mem[16'h1568] <= 0;
        weight_mem[16'h1569] <= 0;
        weight_mem[16'h156A] <= 0;
        weight_mem[16'h156B] <= 0;
        weight_mem[16'h156C] <= 0;
        weight_mem[16'h156D] <= 0;
        weight_mem[16'h156E] <= 0;
        weight_mem[16'h156F] <= 0;
        weight_mem[16'h1570] <= 0;
        weight_mem[16'h1571] <= 0;
        weight_mem[16'h1572] <= 0;
        weight_mem[16'h1573] <= 0;
        weight_mem[16'h1574] <= 0;
        weight_mem[16'h1575] <= 0;
        weight_mem[16'h1576] <= 0;
        weight_mem[16'h1577] <= 0;
        weight_mem[16'h1578] <= 0;
        weight_mem[16'h1579] <= 0;
        weight_mem[16'h157A] <= 0;
        weight_mem[16'h157B] <= 0;
        weight_mem[16'h157C] <= 0;
        weight_mem[16'h157D] <= 0;
        weight_mem[16'h157E] <= 0;
        weight_mem[16'h157F] <= 0;
        weight_mem[16'h1580] <= 0;
        weight_mem[16'h1581] <= 0;
        weight_mem[16'h1582] <= 0;
        weight_mem[16'h1583] <= 0;
        weight_mem[16'h1584] <= 0;
        weight_mem[16'h1585] <= 0;
        weight_mem[16'h1586] <= 0;
        weight_mem[16'h1587] <= 0;
        weight_mem[16'h1588] <= 0;
        weight_mem[16'h1589] <= 0;
        weight_mem[16'h158A] <= 0;
        weight_mem[16'h158B] <= 0;
        weight_mem[16'h158C] <= 0;
        weight_mem[16'h158D] <= 0;
        weight_mem[16'h158E] <= 0;
        weight_mem[16'h158F] <= 0;
        weight_mem[16'h1590] <= 0;
        weight_mem[16'h1591] <= 0;
        weight_mem[16'h1592] <= 0;
        weight_mem[16'h1593] <= 0;
        weight_mem[16'h1594] <= 0;
        weight_mem[16'h1595] <= 0;
        weight_mem[16'h1596] <= 0;
        weight_mem[16'h1597] <= 0;
        weight_mem[16'h1598] <= 0;
        weight_mem[16'h1599] <= 0;
        weight_mem[16'h159A] <= 0;
        weight_mem[16'h159B] <= 0;
        weight_mem[16'h159C] <= 0;
        weight_mem[16'h159D] <= 0;
        weight_mem[16'h159E] <= 0;
        weight_mem[16'h159F] <= 0;
        weight_mem[16'h15A0] <= 0;
        weight_mem[16'h15A1] <= 0;
        weight_mem[16'h15A2] <= 0;
        weight_mem[16'h15A3] <= 0;
        weight_mem[16'h15A4] <= 0;
        weight_mem[16'h15A5] <= 0;
        weight_mem[16'h15A6] <= 0;
        weight_mem[16'h15A7] <= 0;
        weight_mem[16'h15A8] <= 0;
        weight_mem[16'h15A9] <= 0;
        weight_mem[16'h15AA] <= 0;
        weight_mem[16'h15AB] <= 0;
        weight_mem[16'h15AC] <= 0;
        weight_mem[16'h15AD] <= 0;
        weight_mem[16'h15AE] <= 0;
        weight_mem[16'h15AF] <= 0;

        // layer 1 neuron 11
        weight_mem[16'h1600] <= 241;
        weight_mem[16'h1601] <= 241;
        weight_mem[16'h1602] <= 4;
        weight_mem[16'h1603] <= 246;
        weight_mem[16'h1604] <= 5;
        weight_mem[16'h1605] <= 241;
        weight_mem[16'h1606] <= 3;
        weight_mem[16'h1607] <= 237;
        weight_mem[16'h1608] <= 247;
        weight_mem[16'h1609] <= 241;
        weight_mem[16'h160A] <= 254;
        weight_mem[16'h160B] <= 6;
        weight_mem[16'h160C] <= 237;
        weight_mem[16'h160D] <= 8;
        weight_mem[16'h160E] <= 1;
        weight_mem[16'h160F] <= 249;
        weight_mem[16'h1610] <= 3;
        weight_mem[16'h1611] <= 0;
        weight_mem[16'h1612] <= 237;
        weight_mem[16'h1613] <= 2;
        weight_mem[16'h1614] <= 242;
        weight_mem[16'h1615] <= 3;
        weight_mem[16'h1616] <= 238;
        weight_mem[16'h1617] <= 248;
        weight_mem[16'h1618] <= 5;
        weight_mem[16'h1619] <= 247;
        weight_mem[16'h161A] <= 245;
        weight_mem[16'h161B] <= 249;
        weight_mem[16'h161C] <= 244;
        weight_mem[16'h161D] <= 234;
        weight_mem[16'h161E] <= 243;
        weight_mem[16'h161F] <= 254;
        weight_mem[16'h1620] <= 238;
        weight_mem[16'h1621] <= 239;
        weight_mem[16'h1622] <= 230;
        weight_mem[16'h1623] <= 222;
        weight_mem[16'h1624] <= 235;
        weight_mem[16'h1625] <= 236;
        weight_mem[16'h1626] <= 237;
        weight_mem[16'h1627] <= 223;
        weight_mem[16'h1628] <= 234;
        weight_mem[16'h1629] <= 253;
        weight_mem[16'h162A] <= 229;
        weight_mem[16'h162B] <= 246;
        weight_mem[16'h162C] <= 1;
        weight_mem[16'h162D] <= 239;
        weight_mem[16'h162E] <= 255;
        weight_mem[16'h162F] <= 7;
        weight_mem[16'h1630] <= 8;
        weight_mem[16'h1631] <= 254;
        weight_mem[16'h1632] <= 250;
        weight_mem[16'h1633] <= 243;
        weight_mem[16'h1634] <= 253;
        weight_mem[16'h1635] <= 1;
        weight_mem[16'h1636] <= 241;
        weight_mem[16'h1637] <= 230;
        weight_mem[16'h1638] <= 211;
        weight_mem[16'h1639] <= 205;
        weight_mem[16'h163A] <= 233;
        weight_mem[16'h163B] <= 216;
        weight_mem[16'h163C] <= 243;
        weight_mem[16'h163D] <= 253;
        weight_mem[16'h163E] <= 234;
        weight_mem[16'h163F] <= 248;
        weight_mem[16'h1640] <= 229;
        weight_mem[16'h1641] <= 240;
        weight_mem[16'h1642] <= 232;
        weight_mem[16'h1643] <= 235;
        weight_mem[16'h1644] <= 241;
        weight_mem[16'h1645] <= 242;
        weight_mem[16'h1646] <= 242;
        weight_mem[16'h1647] <= 251;
        weight_mem[16'h1648] <= 245;
        weight_mem[16'h1649] <= 247;
        weight_mem[16'h164A] <= 2;
        weight_mem[16'h164B] <= 8;
        weight_mem[16'h164C] <= 2;
        weight_mem[16'h164D] <= 255;
        weight_mem[16'h164E] <= 249;
        weight_mem[16'h164F] <= 242;
        weight_mem[16'h1650] <= 241;
        weight_mem[16'h1651] <= 5;
        weight_mem[16'h1652] <= 3;
        weight_mem[16'h1653] <= 254;
        weight_mem[16'h1654] <= 244;
        weight_mem[16'h1655] <= 241;
        weight_mem[16'h1656] <= 2;
        weight_mem[16'h1657] <= 253;
        weight_mem[16'h1658] <= 11;
        weight_mem[16'h1659] <= 27;
        weight_mem[16'h165A] <= 17;
        weight_mem[16'h165B] <= 10;
        weight_mem[16'h165C] <= 4;
        weight_mem[16'h165D] <= 243;
        weight_mem[16'h165E] <= 8;
        weight_mem[16'h165F] <= 6;
        weight_mem[16'h1660] <= 8;
        weight_mem[16'h1661] <= 3;
        weight_mem[16'h1662] <= 10;
        weight_mem[16'h1663] <= 4;
        weight_mem[16'h1664] <= 6;
        weight_mem[16'h1665] <= 15;
        weight_mem[16'h1666] <= 34;
        weight_mem[16'h1667] <= 39;
        weight_mem[16'h1668] <= 49;
        weight_mem[16'h1669] <= 43;
        weight_mem[16'h166A] <= 42;
        weight_mem[16'h166B] <= 20;
        weight_mem[16'h166C] <= 254;
        weight_mem[16'h166D] <= 13;
        weight_mem[16'h166E] <= 25;
        weight_mem[16'h166F] <= 55;
        weight_mem[16'h1670] <= 83;
        weight_mem[16'h1671] <= 73;
        weight_mem[16'h1672] <= 71;
        weight_mem[16'h1673] <= 51;
        weight_mem[16'h1674] <= 12;
        weight_mem[16'h1675] <= 13;
        weight_mem[16'h1676] <= 1;
        weight_mem[16'h1677] <= 253;
        weight_mem[16'h1678] <= 2;
        weight_mem[16'h1679] <= 249;
        weight_mem[16'h167A] <= 251;
        weight_mem[16'h167B] <= 2;
        weight_mem[16'h167C] <= 25;
        weight_mem[16'h167D] <= 41;
        weight_mem[16'h167E] <= 38;
        weight_mem[16'h167F] <= 49;
        weight_mem[16'h1680] <= 44;
        weight_mem[16'h1681] <= 25;
        weight_mem[16'h1682] <= 29;
        weight_mem[16'h1683] <= 29;
        weight_mem[16'h1684] <= 239;
        weight_mem[16'h1685] <= 9;
        weight_mem[16'h1686] <= 49;
        weight_mem[16'h1687] <= 88;
        weight_mem[16'h1688] <= 109;
        weight_mem[16'h1689] <= 98;
        weight_mem[16'h168A] <= 75;
        weight_mem[16'h168B] <= 70;
        weight_mem[16'h168C] <= 37;
        weight_mem[16'h168D] <= 10;
        weight_mem[16'h168E] <= 244;
        weight_mem[16'h168F] <= 253;
        weight_mem[16'h1690] <= 236;
        weight_mem[16'h1691] <= 3;
        weight_mem[16'h1692] <= 8;
        weight_mem[16'h1693] <= 19;
        weight_mem[16'h1694] <= 19;
        weight_mem[16'h1695] <= 20;
        weight_mem[16'h1696] <= 20;
        weight_mem[16'h1697] <= 2;
        weight_mem[16'h1698] <= 2;
        weight_mem[16'h1699] <= 2;
        weight_mem[16'h169A] <= 11;
        weight_mem[16'h169B] <= 11;
        weight_mem[16'h169C] <= 228;
        weight_mem[16'h169D] <= 27;
        weight_mem[16'h169E] <= 88;
        weight_mem[16'h169F] <= 88;
        weight_mem[16'h16A0] <= 107;
        weight_mem[16'h16A1] <= 84;
        weight_mem[16'h16A2] <= 53;
        weight_mem[16'h16A3] <= 32;
        weight_mem[16'h16A4] <= 20;
        weight_mem[16'h16A5] <= 3;
        weight_mem[16'h16A6] <= 254;
        weight_mem[16'h16A7] <= 241;
        weight_mem[16'h16A8] <= 253;
        weight_mem[16'h16A9] <= 236;
        weight_mem[16'h16AA] <= 255;
        weight_mem[16'h16AB] <= 4;
        weight_mem[16'h16AC] <= 5;
        weight_mem[16'h16AD] <= 4;
        weight_mem[16'h16AE] <= 16;
        weight_mem[16'h16AF] <= 22;
        weight_mem[16'h16B0] <= 16;
        weight_mem[16'h16B1] <= 64;
        weight_mem[16'h16B2] <= 71;
        weight_mem[16'h16B3] <= 39;
        weight_mem[16'h16B4] <= 25;
        weight_mem[16'h16B5] <= 79;
        weight_mem[16'h16B6] <= 77;
        weight_mem[16'h16B7] <= 69;
        weight_mem[16'h16B8] <= 50;
        weight_mem[16'h16B9] <= 34;
        weight_mem[16'h16BA] <= 19;
        weight_mem[16'h16BB] <= 7;
        weight_mem[16'h16BC] <= 0;
        weight_mem[16'h16BD] <= 255;
        weight_mem[16'h16BE] <= 11;
        weight_mem[16'h16BF] <= 244;
        weight_mem[16'h16C0] <= 236;
        weight_mem[16'h16C1] <= 253;
        weight_mem[16'h16C2] <= 247;
        weight_mem[16'h16C3] <= 7;
        weight_mem[16'h16C4] <= 29;
        weight_mem[16'h16C5] <= 17;
        weight_mem[16'h16C6] <= 12;
        weight_mem[16'h16C7] <= 9;
        weight_mem[16'h16C8] <= 6;
        weight_mem[16'h16C9] <= 47;
        weight_mem[16'h16CA] <= 46;
        weight_mem[16'h16CB] <= 255;
        weight_mem[16'h16CC] <= 225;
        weight_mem[16'h16CD] <= 34;
        weight_mem[16'h16CE] <= 55;
        weight_mem[16'h16CF] <= 23;
        weight_mem[16'h16D0] <= 7;
        weight_mem[16'h16D1] <= 255;
        weight_mem[16'h16D2] <= 6;
        weight_mem[16'h16D3] <= 240;
        weight_mem[16'h16D4] <= 239;
        weight_mem[16'h16D5] <= 241;
        weight_mem[16'h16D6] <= 240;
        weight_mem[16'h16D7] <= 238;
        weight_mem[16'h16D8] <= 246;
        weight_mem[16'h16D9] <= 246;
        weight_mem[16'h16DA] <= 3;
        weight_mem[16'h16DB] <= 3;
        weight_mem[16'h16DC] <= 36;
        weight_mem[16'h16DD] <= 17;
        weight_mem[16'h16DE] <= 15;
        weight_mem[16'h16DF] <= 241;
        weight_mem[16'h16E0] <= 216;
        weight_mem[16'h16E1] <= 239;
        weight_mem[16'h16E2] <= 241;
        weight_mem[16'h16E3] <= 205;
        weight_mem[16'h16E4] <= 157;
        weight_mem[16'h16E5] <= 3;
        weight_mem[16'h16E6] <= 59;
        weight_mem[16'h16E7] <= 56;
        weight_mem[16'h16E8] <= 39;
        weight_mem[16'h16E9] <= 11;
        weight_mem[16'h16EA] <= 0;
        weight_mem[16'h16EB] <= 236;
        weight_mem[16'h16EC] <= 228;
        weight_mem[16'h16ED] <= 226;
        weight_mem[16'h16EE] <= 251;
        weight_mem[16'h16EF] <= 253;
        weight_mem[16'h16F0] <= 239;
        weight_mem[16'h16F1] <= 236;
        weight_mem[16'h16F2] <= 8;
        weight_mem[16'h16F3] <= 2;
        weight_mem[16'h16F4] <= 27;
        weight_mem[16'h16F5] <= 11;
        weight_mem[16'h16F6] <= 32;
        weight_mem[16'h16F7] <= 10;
        weight_mem[16'h16F8] <= 216;
        weight_mem[16'h16F9] <= 185;
        weight_mem[16'h16FA] <= 239;
        weight_mem[16'h16FB] <= 203;
        weight_mem[16'h16FC] <= 195;
        weight_mem[16'h16FD] <= 59;
        weight_mem[16'h16FE] <= 90;
        weight_mem[16'h16FF] <= 76;
        weight_mem[16'h1700] <= 1;
        weight_mem[16'h1701] <= 8;
        weight_mem[16'h1702] <= 2;
        weight_mem[16'h1703] <= 236;
        weight_mem[16'h1704] <= 238;
        weight_mem[16'h1705] <= 225;
        weight_mem[16'h1706] <= 250;
        weight_mem[16'h1707] <= 240;
        weight_mem[16'h1708] <= 5;
        weight_mem[16'h1709] <= 246;
        weight_mem[16'h170A] <= 13;
        weight_mem[16'h170B] <= 7;
        weight_mem[16'h170C] <= 13;
        weight_mem[16'h170D] <= 18;
        weight_mem[16'h170E] <= 32;
        weight_mem[16'h170F] <= 245;
        weight_mem[16'h1710] <= 238;
        weight_mem[16'h1711] <= 203;
        weight_mem[16'h1712] <= 240;
        weight_mem[16'h1713] <= 7;
        weight_mem[16'h1714] <= 2;
        weight_mem[16'h1715] <= 35;
        weight_mem[16'h1716] <= 27;
        weight_mem[16'h1717] <= 1;
        weight_mem[16'h1718] <= 231;
        weight_mem[16'h1719] <= 244;
        weight_mem[16'h171A] <= 15;
        weight_mem[16'h171B] <= 254;
        weight_mem[16'h171C] <= 215;
        weight_mem[16'h171D] <= 238;
        weight_mem[16'h171E] <= 235;
        weight_mem[16'h171F] <= 4;
        weight_mem[16'h1720] <= 239;
        weight_mem[16'h1721] <= 250;
        weight_mem[16'h1722] <= 248;
        weight_mem[16'h1723] <= 21;
        weight_mem[16'h1724] <= 22;
        weight_mem[16'h1725] <= 46;
        weight_mem[16'h1726] <= 14;
        weight_mem[16'h1727] <= 2;
        weight_mem[16'h1728] <= 230;
        weight_mem[16'h1729] <= 184;
        weight_mem[16'h172A] <= 166;
        weight_mem[16'h172B] <= 185;
        weight_mem[16'h172C] <= 181;
        weight_mem[16'h172D] <= 185;
        weight_mem[16'h172E] <= 182;
        weight_mem[16'h172F] <= 185;
        weight_mem[16'h1730] <= 225;
        weight_mem[16'h1731] <= 219;
        weight_mem[16'h1732] <= 239;
        weight_mem[16'h1733] <= 242;
        weight_mem[16'h1734] <= 229;
        weight_mem[16'h1735] <= 242;
        weight_mem[16'h1736] <= 237;
        weight_mem[16'h1737] <= 252;
        weight_mem[16'h1738] <= 248;
        weight_mem[16'h1739] <= 252;
        weight_mem[16'h173A] <= 243;
        weight_mem[16'h173B] <= 11;
        weight_mem[16'h173C] <= 7;
        weight_mem[16'h173D] <= 16;
        weight_mem[16'h173E] <= 249;
        weight_mem[16'h173F] <= 254;
        weight_mem[16'h1740] <= 230;
        weight_mem[16'h1741] <= 191;
        weight_mem[16'h1742] <= 171;
        weight_mem[16'h1743] <= 143;
        weight_mem[16'h1744] <= 128;
        weight_mem[16'h1745] <= 150;
        weight_mem[16'h1746] <= 184;
        weight_mem[16'h1747] <= 181;
        weight_mem[16'h1748] <= 190;
        weight_mem[16'h1749] <= 231;
        weight_mem[16'h174A] <= 236;
        weight_mem[16'h174B] <= 228;
        weight_mem[16'h174C] <= 237;
        weight_mem[16'h174D] <= 233;
        weight_mem[16'h174E] <= 0;
        weight_mem[16'h174F] <= 250;
        weight_mem[16'h1750] <= 237;
        weight_mem[16'h1751] <= 236;
        weight_mem[16'h1752] <= 243;
        weight_mem[16'h1753] <= 6;
        weight_mem[16'h1754] <= 246;
        weight_mem[16'h1755] <= 248;
        weight_mem[16'h1756] <= 10;
        weight_mem[16'h1757] <= 246;
        weight_mem[16'h1758] <= 236;
        weight_mem[16'h1759] <= 4;
        weight_mem[16'h175A] <= 10;
        weight_mem[16'h175B] <= 20;
        weight_mem[16'h175C] <= 10;
        weight_mem[16'h175D] <= 17;
        weight_mem[16'h175E] <= 13;
        weight_mem[16'h175F] <= 242;
        weight_mem[16'h1760] <= 234;
        weight_mem[16'h1761] <= 245;
        weight_mem[16'h1762] <= 246;
        weight_mem[16'h1763] <= 240;
        weight_mem[16'h1764] <= 242;
        weight_mem[16'h1765] <= 235;
        weight_mem[16'h1766] <= 5;
        weight_mem[16'h1767] <= 0;
        weight_mem[16'h1768] <= 3;
        weight_mem[16'h1769] <= 249;
        weight_mem[16'h176A] <= 6;
        weight_mem[16'h176B] <= 245;
        weight_mem[16'h176C] <= 243;
        weight_mem[16'h176D] <= 15;
        weight_mem[16'h176E] <= 15;
        weight_mem[16'h176F] <= 40;
        weight_mem[16'h1770] <= 37;
        weight_mem[16'h1771] <= 40;
        weight_mem[16'h1772] <= 57;
        weight_mem[16'h1773] <= 78;
        weight_mem[16'h1774] <= 75;
        weight_mem[16'h1775] <= 50;
        weight_mem[16'h1776] <= 53;
        weight_mem[16'h1777] <= 47;
        weight_mem[16'h1778] <= 25;
        weight_mem[16'h1779] <= 6;
        weight_mem[16'h177A] <= 7;
        weight_mem[16'h177B] <= 8;
        weight_mem[16'h177C] <= 246;
        weight_mem[16'h177D] <= 239;
        weight_mem[16'h177E] <= 252;
        weight_mem[16'h177F] <= 243;
        weight_mem[16'h1780] <= 248;
        weight_mem[16'h1781] <= 235;
        weight_mem[16'h1782] <= 7;
        weight_mem[16'h1783] <= 10;
        weight_mem[16'h1784] <= 250;
        weight_mem[16'h1785] <= 5;
        weight_mem[16'h1786] <= 10;
        weight_mem[16'h1787] <= 7;
        weight_mem[16'h1788] <= 13;
        weight_mem[16'h1789] <= 30;
        weight_mem[16'h178A] <= 35;
        weight_mem[16'h178B] <= 45;
        weight_mem[16'h178C] <= 34;
        weight_mem[16'h178D] <= 45;
        weight_mem[16'h178E] <= 33;
        weight_mem[16'h178F] <= 32;
        weight_mem[16'h1790] <= 22;
        weight_mem[16'h1791] <= 9;
        weight_mem[16'h1792] <= 247;
        weight_mem[16'h1793] <= 3;
        weight_mem[16'h1794] <= 246;
        weight_mem[16'h1795] <= 236;
        weight_mem[16'h1796] <= 244;
        weight_mem[16'h1797] <= 1;
        weight_mem[16'h1798] <= 249;
        weight_mem[16'h1799] <= 0;
        weight_mem[16'h179A] <= 237;
        weight_mem[16'h179B] <= 250;
        weight_mem[16'h179C] <= 250;
        weight_mem[16'h179D] <= 251;
        weight_mem[16'h179E] <= 247;
        weight_mem[16'h179F] <= 0;
        weight_mem[16'h17A0] <= 11;
        weight_mem[16'h17A1] <= 242;
        weight_mem[16'h17A2] <= 248;
        weight_mem[16'h17A3] <= 0;
        weight_mem[16'h17A4] <= 12;
        weight_mem[16'h17A5] <= 2;
        weight_mem[16'h17A6] <= 242;
        weight_mem[16'h17A7] <= 255;
        weight_mem[16'h17A8] <= 254;
        weight_mem[16'h17A9] <= 245;
        weight_mem[16'h17AA] <= 9;
        weight_mem[16'h17AB] <= 236;
        weight_mem[16'h17AC] <= 247;
        weight_mem[16'h17AD] <= 4;
        weight_mem[16'h17AE] <= 250;
        weight_mem[16'h17AF] <= 1;

        // layer 1 neuron 12
        weight_mem[16'h1800] <= 176;
        weight_mem[16'h1801] <= 176;
        weight_mem[16'h1802] <= 176;
        weight_mem[16'h1803] <= 176;
        weight_mem[16'h1804] <= 176;
        weight_mem[16'h1805] <= 176;
        weight_mem[16'h1806] <= 176;
        weight_mem[16'h1807] <= 176;
        weight_mem[16'h1808] <= 176;
        weight_mem[16'h1809] <= 176;
        weight_mem[16'h180A] <= 176;
        weight_mem[16'h180B] <= 176;
        weight_mem[16'h180C] <= 176;
        weight_mem[16'h180D] <= 176;
        weight_mem[16'h180E] <= 176;
        weight_mem[16'h180F] <= 176;
        weight_mem[16'h1810] <= 176;
        weight_mem[16'h1811] <= 176;
        weight_mem[16'h1812] <= 176;
        weight_mem[16'h1813] <= 176;
        weight_mem[16'h1814] <= 176;
        weight_mem[16'h1815] <= 176;
        weight_mem[16'h1816] <= 176;
        weight_mem[16'h1817] <= 176;
        weight_mem[16'h1818] <= 176;
        weight_mem[16'h1819] <= 176;
        weight_mem[16'h181A] <= 176;
        weight_mem[16'h181B] <= 176;
        weight_mem[16'h181C] <= 176;
        weight_mem[16'h181D] <= 176;
        weight_mem[16'h181E] <= 176;
        weight_mem[16'h181F] <= 176;
        weight_mem[16'h1820] <= 176;
        weight_mem[16'h1821] <= 176;
        weight_mem[16'h1822] <= 178;
        weight_mem[16'h1823] <= 179;
        weight_mem[16'h1824] <= 178;
        weight_mem[16'h1825] <= 178;
        weight_mem[16'h1826] <= 178;
        weight_mem[16'h1827] <= 179;
        weight_mem[16'h1828] <= 178;
        weight_mem[16'h1829] <= 178;
        weight_mem[16'h182A] <= 179;
        weight_mem[16'h182B] <= 178;
        weight_mem[16'h182C] <= 176;
        weight_mem[16'h182D] <= 176;
        weight_mem[16'h182E] <= 176;
        weight_mem[16'h182F] <= 176;
        weight_mem[16'h1830] <= 176;
        weight_mem[16'h1831] <= 176;
        weight_mem[16'h1832] <= 176;
        weight_mem[16'h1833] <= 176;
        weight_mem[16'h1834] <= 177;
        weight_mem[16'h1835] <= 177;
        weight_mem[16'h1836] <= 177;
        weight_mem[16'h1837] <= 178;
        weight_mem[16'h1838] <= 176;
        weight_mem[16'h1839] <= 177;
        weight_mem[16'h183A] <= 182;
        weight_mem[16'h183B] <= 189;
        weight_mem[16'h183C] <= 193;
        weight_mem[16'h183D] <= 186;
        weight_mem[16'h183E] <= 186;
        weight_mem[16'h183F] <= 189;
        weight_mem[16'h1840] <= 185;
        weight_mem[16'h1841] <= 183;
        weight_mem[16'h1842] <= 181;
        weight_mem[16'h1843] <= 178;
        weight_mem[16'h1844] <= 176;
        weight_mem[16'h1845] <= 176;
        weight_mem[16'h1846] <= 176;
        weight_mem[16'h1847] <= 176;
        weight_mem[16'h1848] <= 176;
        weight_mem[16'h1849] <= 176;
        weight_mem[16'h184A] <= 176;
        weight_mem[16'h184B] <= 177;
        weight_mem[16'h184C] <= 178;
        weight_mem[16'h184D] <= 177;
        weight_mem[16'h184E] <= 180;
        weight_mem[16'h184F] <= 184;
        weight_mem[16'h1850] <= 186;
        weight_mem[16'h1851] <= 188;
        weight_mem[16'h1852] <= 199;
        weight_mem[16'h1853] <= 215;
        weight_mem[16'h1854] <= 220;
        weight_mem[16'h1855] <= 212;
        weight_mem[16'h1856] <= 203;
        weight_mem[16'h1857] <= 205;
        weight_mem[16'h1858] <= 213;
        weight_mem[16'h1859] <= 220;
        weight_mem[16'h185A] <= 207;
        weight_mem[16'h185B] <= 186;
        weight_mem[16'h185C] <= 172;
        weight_mem[16'h185D] <= 167;
        weight_mem[16'h185E] <= 168;
        weight_mem[16'h185F] <= 173;
        weight_mem[16'h1860] <= 176;
        weight_mem[16'h1861] <= 176;
        weight_mem[16'h1862] <= 178;
        weight_mem[16'h1863] <= 179;
        weight_mem[16'h1864] <= 179;
        weight_mem[16'h1865] <= 177;
        weight_mem[16'h1866] <= 195;
        weight_mem[16'h1867] <= 205;
        weight_mem[16'h1868] <= 214;
        weight_mem[16'h1869] <= 225;
        weight_mem[16'h186A] <= 240;
        weight_mem[16'h186B] <= 241;
        weight_mem[16'h186C] <= 241;
        weight_mem[16'h186D] <= 225;
        weight_mem[16'h186E] <= 217;
        weight_mem[16'h186F] <= 206;
        weight_mem[16'h1870] <= 218;
        weight_mem[16'h1871] <= 243;
        weight_mem[16'h1872] <= 226;
        weight_mem[16'h1873] <= 193;
        weight_mem[16'h1874] <= 184;
        weight_mem[16'h1875] <= 171;
        weight_mem[16'h1876] <= 158;
        weight_mem[16'h1877] <= 163;
        weight_mem[16'h1878] <= 176;
        weight_mem[16'h1879] <= 176;
        weight_mem[16'h187A] <= 179;
        weight_mem[16'h187B] <= 183;
        weight_mem[16'h187C] <= 187;
        weight_mem[16'h187D] <= 187;
        weight_mem[16'h187E] <= 202;
        weight_mem[16'h187F] <= 198;
        weight_mem[16'h1880] <= 213;
        weight_mem[16'h1881] <= 236;
        weight_mem[16'h1882] <= 238;
        weight_mem[16'h1883] <= 226;
        weight_mem[16'h1884] <= 206;
        weight_mem[16'h1885] <= 197;
        weight_mem[16'h1886] <= 214;
        weight_mem[16'h1887] <= 231;
        weight_mem[16'h1888] <= 221;
        weight_mem[16'h1889] <= 213;
        weight_mem[16'h188A] <= 184;
        weight_mem[16'h188B] <= 179;
        weight_mem[16'h188C] <= 184;
        weight_mem[16'h188D] <= 186;
        weight_mem[16'h188E] <= 177;
        weight_mem[16'h188F] <= 175;
        weight_mem[16'h1890] <= 176;
        weight_mem[16'h1891] <= 177;
        weight_mem[16'h1892] <= 180;
        weight_mem[16'h1893] <= 185;
        weight_mem[16'h1894] <= 192;
        weight_mem[16'h1895] <= 187;
        weight_mem[16'h1896] <= 183;
        weight_mem[16'h1897] <= 180;
        weight_mem[16'h1898] <= 214;
        weight_mem[16'h1899] <= 242;
        weight_mem[16'h189A] <= 240;
        weight_mem[16'h189B] <= 238;
        weight_mem[16'h189C] <= 230;
        weight_mem[16'h189D] <= 221;
        weight_mem[16'h189E] <= 232;
        weight_mem[16'h189F] <= 250;
        weight_mem[16'h18A0] <= 240;
        weight_mem[16'h18A1] <= 208;
        weight_mem[16'h18A2] <= 176;
        weight_mem[16'h18A3] <= 183;
        weight_mem[16'h18A4] <= 181;
        weight_mem[16'h18A5] <= 183;
        weight_mem[16'h18A6] <= 181;
        weight_mem[16'h18A7] <= 178;
        weight_mem[16'h18A8] <= 176;
        weight_mem[16'h18A9] <= 177;
        weight_mem[16'h18AA] <= 178;
        weight_mem[16'h18AB] <= 187;
        weight_mem[16'h18AC] <= 186;
        weight_mem[16'h18AD] <= 187;
        weight_mem[16'h18AE] <= 206;
        weight_mem[16'h18AF] <= 214;
        weight_mem[16'h18B0] <= 237;
        weight_mem[16'h18B1] <= 250;
        weight_mem[16'h18B2] <= 250;
        weight_mem[16'h18B3] <= 243;
        weight_mem[16'h18B4] <= 238;
        weight_mem[16'h18B5] <= 241;
        weight_mem[16'h18B6] <= 246;
        weight_mem[16'h18B7] <= 247;
        weight_mem[16'h18B8] <= 234;
        weight_mem[16'h18B9] <= 194;
        weight_mem[16'h18BA] <= 178;
        weight_mem[16'h18BB] <= 185;
        weight_mem[16'h18BC] <= 184;
        weight_mem[16'h18BD] <= 184;
        weight_mem[16'h18BE] <= 180;
        weight_mem[16'h18BF] <= 177;
        weight_mem[16'h18C0] <= 176;
        weight_mem[16'h18C1] <= 176;
        weight_mem[16'h18C2] <= 177;
        weight_mem[16'h18C3] <= 185;
        weight_mem[16'h18C4] <= 186;
        weight_mem[16'h18C5] <= 188;
        weight_mem[16'h18C6] <= 220;
        weight_mem[16'h18C7] <= 222;
        weight_mem[16'h18C8] <= 213;
        weight_mem[16'h18C9] <= 211;
        weight_mem[16'h18CA] <= 222;
        weight_mem[16'h18CB] <= 222;
        weight_mem[16'h18CC] <= 244;
        weight_mem[16'h18CD] <= 249;
        weight_mem[16'h18CE] <= 245;
        weight_mem[16'h18CF] <= 237;
        weight_mem[16'h18D0] <= 219;
        weight_mem[16'h18D1] <= 181;
        weight_mem[16'h18D2] <= 164;
        weight_mem[16'h18D3] <= 169;
        weight_mem[16'h18D4] <= 175;
        weight_mem[16'h18D5] <= 176;
        weight_mem[16'h18D6] <= 177;
        weight_mem[16'h18D7] <= 176;
        weight_mem[16'h18D8] <= 176;
        weight_mem[16'h18D9] <= 176;
        weight_mem[16'h18DA] <= 176;
        weight_mem[16'h18DB] <= 184;
        weight_mem[16'h18DC] <= 187;
        weight_mem[16'h18DD] <= 192;
        weight_mem[16'h18DE] <= 210;
        weight_mem[16'h18DF] <= 212;
        weight_mem[16'h18E0] <= 173;
        weight_mem[16'h18E1] <= 128;
        weight_mem[16'h18E2] <= 161;
        weight_mem[16'h18E3] <= 193;
        weight_mem[16'h18E4] <= 219;
        weight_mem[16'h18E5] <= 235;
        weight_mem[16'h18E6] <= 237;
        weight_mem[16'h18E7] <= 238;
        weight_mem[16'h18E8] <= 215;
        weight_mem[16'h18E9] <= 190;
        weight_mem[16'h18EA] <= 171;
        weight_mem[16'h18EB] <= 168;
        weight_mem[16'h18EC] <= 172;
        weight_mem[16'h18ED] <= 174;
        weight_mem[16'h18EE] <= 176;
        weight_mem[16'h18EF] <= 176;
        weight_mem[16'h18F0] <= 176;
        weight_mem[16'h18F1] <= 176;
        weight_mem[16'h18F2] <= 176;
        weight_mem[16'h18F3] <= 183;
        weight_mem[16'h18F4] <= 190;
        weight_mem[16'h18F5] <= 201;
        weight_mem[16'h18F6] <= 200;
        weight_mem[16'h18F7] <= 193;
        weight_mem[16'h18F8] <= 158;
        weight_mem[16'h18F9] <= 152;
        weight_mem[16'h18FA] <= 179;
        weight_mem[16'h18FB] <= 201;
        weight_mem[16'h18FC] <= 208;
        weight_mem[16'h18FD] <= 212;
        weight_mem[16'h18FE] <= 221;
        weight_mem[16'h18FF] <= 234;
        weight_mem[16'h1900] <= 222;
        weight_mem[16'h1901] <= 213;
        weight_mem[16'h1902] <= 197;
        weight_mem[16'h1903] <= 188;
        weight_mem[16'h1904] <= 179;
        weight_mem[16'h1905] <= 173;
        weight_mem[16'h1906] <= 176;
        weight_mem[16'h1907] <= 176;
        weight_mem[16'h1908] <= 176;
        weight_mem[16'h1909] <= 176;
        weight_mem[16'h190A] <= 175;
        weight_mem[16'h190B] <= 186;
        weight_mem[16'h190C] <= 194;
        weight_mem[16'h190D] <= 194;
        weight_mem[16'h190E] <= 198;
        weight_mem[16'h190F] <= 200;
        weight_mem[16'h1910] <= 188;
        weight_mem[16'h1911] <= 202;
        weight_mem[16'h1912] <= 212;
        weight_mem[16'h1913] <= 201;
        weight_mem[16'h1914] <= 202;
        weight_mem[16'h1915] <= 227;
        weight_mem[16'h1916] <= 223;
        weight_mem[16'h1917] <= 225;
        weight_mem[16'h1918] <= 221;
        weight_mem[16'h1919] <= 219;
        weight_mem[16'h191A] <= 211;
        weight_mem[16'h191B] <= 193;
        weight_mem[16'h191C] <= 179;
        weight_mem[16'h191D] <= 174;
        weight_mem[16'h191E] <= 176;
        weight_mem[16'h191F] <= 176;
        weight_mem[16'h1920] <= 176;
        weight_mem[16'h1921] <= 176;
        weight_mem[16'h1922] <= 175;
        weight_mem[16'h1923] <= 189;
        weight_mem[16'h1924] <= 203;
        weight_mem[16'h1925] <= 201;
        weight_mem[16'h1926] <= 206;
        weight_mem[16'h1927] <= 202;
        weight_mem[16'h1928] <= 202;
        weight_mem[16'h1929] <= 219;
        weight_mem[16'h192A] <= 219;
        weight_mem[16'h192B] <= 211;
        weight_mem[16'h192C] <= 239;
        weight_mem[16'h192D] <= 249;
        weight_mem[16'h192E] <= 235;
        weight_mem[16'h192F] <= 216;
        weight_mem[16'h1930] <= 200;
        weight_mem[16'h1931] <= 211;
        weight_mem[16'h1932] <= 208;
        weight_mem[16'h1933] <= 191;
        weight_mem[16'h1934] <= 177;
        weight_mem[16'h1935] <= 175;
        weight_mem[16'h1936] <= 176;
        weight_mem[16'h1937] <= 176;
        weight_mem[16'h1938] <= 176;
        weight_mem[16'h1939] <= 176;
        weight_mem[16'h193A] <= 175;
        weight_mem[16'h193B] <= 181;
        weight_mem[16'h193C] <= 194;
        weight_mem[16'h193D] <= 203;
        weight_mem[16'h193E] <= 216;
        weight_mem[16'h193F] <= 222;
        weight_mem[16'h1940] <= 228;
        weight_mem[16'h1941] <= 211;
        weight_mem[16'h1942] <= 196;
        weight_mem[16'h1943] <= 222;
        weight_mem[16'h1944] <= 244;
        weight_mem[16'h1945] <= 244;
        weight_mem[16'h1946] <= 236;
        weight_mem[16'h1947] <= 223;
        weight_mem[16'h1948] <= 197;
        weight_mem[16'h1949] <= 183;
        weight_mem[16'h194A] <= 195;
        weight_mem[16'h194B] <= 188;
        weight_mem[16'h194C] <= 178;
        weight_mem[16'h194D] <= 175;
        weight_mem[16'h194E] <= 175;
        weight_mem[16'h194F] <= 176;
        weight_mem[16'h1950] <= 176;
        weight_mem[16'h1951] <= 176;
        weight_mem[16'h1952] <= 176;
        weight_mem[16'h1953] <= 176;
        weight_mem[16'h1954] <= 179;
        weight_mem[16'h1955] <= 192;
        weight_mem[16'h1956] <= 210;
        weight_mem[16'h1957] <= 217;
        weight_mem[16'h1958] <= 217;
        weight_mem[16'h1959] <= 196;
        weight_mem[16'h195A] <= 193;
        weight_mem[16'h195B] <= 197;
        weight_mem[16'h195C] <= 210;
        weight_mem[16'h195D] <= 203;
        weight_mem[16'h195E] <= 217;
        weight_mem[16'h195F] <= 218;
        weight_mem[16'h1960] <= 187;
        weight_mem[16'h1961] <= 167;
        weight_mem[16'h1962] <= 183;
        weight_mem[16'h1963] <= 180;
        weight_mem[16'h1964] <= 176;
        weight_mem[16'h1965] <= 176;
        weight_mem[16'h1966] <= 176;
        weight_mem[16'h1967] <= 176;
        weight_mem[16'h1968] <= 176;
        weight_mem[16'h1969] <= 176;
        weight_mem[16'h196A] <= 176;
        weight_mem[16'h196B] <= 176;
        weight_mem[16'h196C] <= 181;
        weight_mem[16'h196D] <= 195;
        weight_mem[16'h196E] <= 201;
        weight_mem[16'h196F] <= 200;
        weight_mem[16'h1970] <= 188;
        weight_mem[16'h1971] <= 193;
        weight_mem[16'h1972] <= 201;
        weight_mem[16'h1973] <= 173;
        weight_mem[16'h1974] <= 142;
        weight_mem[16'h1975] <= 138;
        weight_mem[16'h1976] <= 169;
        weight_mem[16'h1977] <= 192;
        weight_mem[16'h1978] <= 184;
        weight_mem[16'h1979] <= 181;
        weight_mem[16'h197A] <= 182;
        weight_mem[16'h197B] <= 176;
        weight_mem[16'h197C] <= 176;
        weight_mem[16'h197D] <= 176;
        weight_mem[16'h197E] <= 176;
        weight_mem[16'h197F] <= 176;
        weight_mem[16'h1980] <= 176;
        weight_mem[16'h1981] <= 176;
        weight_mem[16'h1982] <= 176;
        weight_mem[16'h1983] <= 176;
        weight_mem[16'h1984] <= 181;
        weight_mem[16'h1985] <= 194;
        weight_mem[16'h1986] <= 193;
        weight_mem[16'h1987] <= 184;
        weight_mem[16'h1988] <= 184;
        weight_mem[16'h1989] <= 194;
        weight_mem[16'h198A] <= 208;
        weight_mem[16'h198B] <= 201;
        weight_mem[16'h198C] <= 168;
        weight_mem[16'h198D] <= 151;
        weight_mem[16'h198E] <= 163;
        weight_mem[16'h198F] <= 185;
        weight_mem[16'h1990] <= 189;
        weight_mem[16'h1991] <= 185;
        weight_mem[16'h1992] <= 180;
        weight_mem[16'h1993] <= 176;
        weight_mem[16'h1994] <= 176;
        weight_mem[16'h1995] <= 176;
        weight_mem[16'h1996] <= 176;
        weight_mem[16'h1997] <= 176;
        weight_mem[16'h1998] <= 176;
        weight_mem[16'h1999] <= 176;
        weight_mem[16'h199A] <= 176;
        weight_mem[16'h199B] <= 176;
        weight_mem[16'h199C] <= 176;
        weight_mem[16'h199D] <= 177;
        weight_mem[16'h199E] <= 177;
        weight_mem[16'h199F] <= 176;
        weight_mem[16'h19A0] <= 178;
        weight_mem[16'h19A1] <= 181;
        weight_mem[16'h19A2] <= 181;
        weight_mem[16'h19A3] <= 179;
        weight_mem[16'h19A4] <= 178;
        weight_mem[16'h19A5] <= 180;
        weight_mem[16'h19A6] <= 182;
        weight_mem[16'h19A7] <= 182;
        weight_mem[16'h19A8] <= 179;
        weight_mem[16'h19A9] <= 176;
        weight_mem[16'h19AA] <= 176;
        weight_mem[16'h19AB] <= 176;
        weight_mem[16'h19AC] <= 176;
        weight_mem[16'h19AD] <= 176;
        weight_mem[16'h19AE] <= 176;
        weight_mem[16'h19AF] <= 176;

        // layer 1 neuron 13
        weight_mem[16'h1A00] <= 167;
        weight_mem[16'h1A01] <= 167;
        weight_mem[16'h1A02] <= 167;
        weight_mem[16'h1A03] <= 167;
        weight_mem[16'h1A04] <= 167;
        weight_mem[16'h1A05] <= 167;
        weight_mem[16'h1A06] <= 167;
        weight_mem[16'h1A07] <= 167;
        weight_mem[16'h1A08] <= 167;
        weight_mem[16'h1A09] <= 167;
        weight_mem[16'h1A0A] <= 167;
        weight_mem[16'h1A0B] <= 167;
        weight_mem[16'h1A0C] <= 167;
        weight_mem[16'h1A0D] <= 167;
        weight_mem[16'h1A0E] <= 167;
        weight_mem[16'h1A0F] <= 167;
        weight_mem[16'h1A10] <= 167;
        weight_mem[16'h1A11] <= 167;
        weight_mem[16'h1A12] <= 167;
        weight_mem[16'h1A13] <= 167;
        weight_mem[16'h1A14] <= 167;
        weight_mem[16'h1A15] <= 167;
        weight_mem[16'h1A16] <= 167;
        weight_mem[16'h1A17] <= 167;
        weight_mem[16'h1A18] <= 167;
        weight_mem[16'h1A19] <= 167;
        weight_mem[16'h1A1A] <= 167;
        weight_mem[16'h1A1B] <= 167;
        weight_mem[16'h1A1C] <= 167;
        weight_mem[16'h1A1D] <= 167;
        weight_mem[16'h1A1E] <= 166;
        weight_mem[16'h1A1F] <= 165;
        weight_mem[16'h1A20] <= 166;
        weight_mem[16'h1A21] <= 167;
        weight_mem[16'h1A22] <= 167;
        weight_mem[16'h1A23] <= 165;
        weight_mem[16'h1A24] <= 165;
        weight_mem[16'h1A25] <= 165;
        weight_mem[16'h1A26] <= 163;
        weight_mem[16'h1A27] <= 161;
        weight_mem[16'h1A28] <= 162;
        weight_mem[16'h1A29] <= 166;
        weight_mem[16'h1A2A] <= 167;
        weight_mem[16'h1A2B] <= 167;
        weight_mem[16'h1A2C] <= 167;
        weight_mem[16'h1A2D] <= 167;
        weight_mem[16'h1A2E] <= 167;
        weight_mem[16'h1A2F] <= 167;
        weight_mem[16'h1A30] <= 167;
        weight_mem[16'h1A31] <= 167;
        weight_mem[16'h1A32] <= 167;
        weight_mem[16'h1A33] <= 167;
        weight_mem[16'h1A34] <= 167;
        weight_mem[16'h1A35] <= 167;
        weight_mem[16'h1A36] <= 161;
        weight_mem[16'h1A37] <= 155;
        weight_mem[16'h1A38] <= 161;
        weight_mem[16'h1A39] <= 162;
        weight_mem[16'h1A3A] <= 163;
        weight_mem[16'h1A3B] <= 161;
        weight_mem[16'h1A3C] <= 168;
        weight_mem[16'h1A3D] <= 171;
        weight_mem[16'h1A3E] <= 142;
        weight_mem[16'h1A3F] <= 128;
        weight_mem[16'h1A40] <= 142;
        weight_mem[16'h1A41] <= 164;
        weight_mem[16'h1A42] <= 169;
        weight_mem[16'h1A43] <= 168;
        weight_mem[16'h1A44] <= 168;
        weight_mem[16'h1A45] <= 167;
        weight_mem[16'h1A46] <= 167;
        weight_mem[16'h1A47] <= 167;
        weight_mem[16'h1A48] <= 167;
        weight_mem[16'h1A49] <= 167;
        weight_mem[16'h1A4A] <= 167;
        weight_mem[16'h1A4B] <= 167;
        weight_mem[16'h1A4C] <= 167;
        weight_mem[16'h1A4D] <= 170;
        weight_mem[16'h1A4E] <= 167;
        weight_mem[16'h1A4F] <= 182;
        weight_mem[16'h1A50] <= 211;
        weight_mem[16'h1A51] <= 222;
        weight_mem[16'h1A52] <= 221;
        weight_mem[16'h1A53] <= 230;
        weight_mem[16'h1A54] <= 236;
        weight_mem[16'h1A55] <= 212;
        weight_mem[16'h1A56] <= 204;
        weight_mem[16'h1A57] <= 200;
        weight_mem[16'h1A58] <= 205;
        weight_mem[16'h1A59] <= 210;
        weight_mem[16'h1A5A] <= 202;
        weight_mem[16'h1A5B] <= 192;
        weight_mem[16'h1A5C] <= 178;
        weight_mem[16'h1A5D] <= 169;
        weight_mem[16'h1A5E] <= 167;
        weight_mem[16'h1A5F] <= 167;
        weight_mem[16'h1A60] <= 167;
        weight_mem[16'h1A61] <= 167;
        weight_mem[16'h1A62] <= 167;
        weight_mem[16'h1A63] <= 169;
        weight_mem[16'h1A64] <= 178;
        weight_mem[16'h1A65] <= 190;
        weight_mem[16'h1A66] <= 196;
        weight_mem[16'h1A67] <= 226;
        weight_mem[16'h1A68] <= 242;
        weight_mem[16'h1A69] <= 249;
        weight_mem[16'h1A6A] <= 252;
        weight_mem[16'h1A6B] <= 254;
        weight_mem[16'h1A6C] <= 253;
        weight_mem[16'h1A6D] <= 241;
        weight_mem[16'h1A6E] <= 242;
        weight_mem[16'h1A6F] <= 248;
        weight_mem[16'h1A70] <= 246;
        weight_mem[16'h1A71] <= 234;
        weight_mem[16'h1A72] <= 220;
        weight_mem[16'h1A73] <= 209;
        weight_mem[16'h1A74] <= 190;
        weight_mem[16'h1A75] <= 172;
        weight_mem[16'h1A76] <= 168;
        weight_mem[16'h1A77] <= 167;
        weight_mem[16'h1A78] <= 167;
        weight_mem[16'h1A79] <= 167;
        weight_mem[16'h1A7A] <= 167;
        weight_mem[16'h1A7B] <= 174;
        weight_mem[16'h1A7C] <= 187;
        weight_mem[16'h1A7D] <= 203;
        weight_mem[16'h1A7E] <= 217;
        weight_mem[16'h1A7F] <= 235;
        weight_mem[16'h1A80] <= 239;
        weight_mem[16'h1A81] <= 245;
        weight_mem[16'h1A82] <= 250;
        weight_mem[16'h1A83] <= 248;
        weight_mem[16'h1A84] <= 247;
        weight_mem[16'h1A85] <= 242;
        weight_mem[16'h1A86] <= 235;
        weight_mem[16'h1A87] <= 237;
        weight_mem[16'h1A88] <= 234;
        weight_mem[16'h1A89] <= 212;
        weight_mem[16'h1A8A] <= 209;
        weight_mem[16'h1A8B] <= 211;
        weight_mem[16'h1A8C] <= 194;
        weight_mem[16'h1A8D] <= 170;
        weight_mem[16'h1A8E] <= 168;
        weight_mem[16'h1A8F] <= 167;
        weight_mem[16'h1A90] <= 167;
        weight_mem[16'h1A91] <= 167;
        weight_mem[16'h1A92] <= 169;
        weight_mem[16'h1A93] <= 171;
        weight_mem[16'h1A94] <= 177;
        weight_mem[16'h1A95] <= 195;
        weight_mem[16'h1A96] <= 213;
        weight_mem[16'h1A97] <= 224;
        weight_mem[16'h1A98] <= 226;
        weight_mem[16'h1A99] <= 243;
        weight_mem[16'h1A9A] <= 250;
        weight_mem[16'h1A9B] <= 251;
        weight_mem[16'h1A9C] <= 251;
        weight_mem[16'h1A9D] <= 250;
        weight_mem[16'h1A9E] <= 244;
        weight_mem[16'h1A9F] <= 231;
        weight_mem[16'h1AA0] <= 214;
        weight_mem[16'h1AA1] <= 201;
        weight_mem[16'h1AA2] <= 203;
        weight_mem[16'h1AA3] <= 209;
        weight_mem[16'h1AA4] <= 193;
        weight_mem[16'h1AA5] <= 171;
        weight_mem[16'h1AA6] <= 168;
        weight_mem[16'h1AA7] <= 167;
        weight_mem[16'h1AA8] <= 167;
        weight_mem[16'h1AA9] <= 167;
        weight_mem[16'h1AAA] <= 168;
        weight_mem[16'h1AAB] <= 169;
        weight_mem[16'h1AAC] <= 177;
        weight_mem[16'h1AAD] <= 194;
        weight_mem[16'h1AAE] <= 203;
        weight_mem[16'h1AAF] <= 209;
        weight_mem[16'h1AB0] <= 224;
        weight_mem[16'h1AB1] <= 242;
        weight_mem[16'h1AB2] <= 245;
        weight_mem[16'h1AB3] <= 248;
        weight_mem[16'h1AB4] <= 250;
        weight_mem[16'h1AB5] <= 250;
        weight_mem[16'h1AB6] <= 250;
        weight_mem[16'h1AB7] <= 249;
        weight_mem[16'h1AB8] <= 232;
        weight_mem[16'h1AB9] <= 213;
        weight_mem[16'h1ABA] <= 204;
        weight_mem[16'h1ABB] <= 202;
        weight_mem[16'h1ABC] <= 183;
        weight_mem[16'h1ABD] <= 169;
        weight_mem[16'h1ABE] <= 168;
        weight_mem[16'h1ABF] <= 167;
        weight_mem[16'h1AC0] <= 167;
        weight_mem[16'h1AC1] <= 167;
        weight_mem[16'h1AC2] <= 162;
        weight_mem[16'h1AC3] <= 163;
        weight_mem[16'h1AC4] <= 182;
        weight_mem[16'h1AC5] <= 199;
        weight_mem[16'h1AC6] <= 198;
        weight_mem[16'h1AC7] <= 199;
        weight_mem[16'h1AC8] <= 233;
        weight_mem[16'h1AC9] <= 246;
        weight_mem[16'h1ACA] <= 244;
        weight_mem[16'h1ACB] <= 248;
        weight_mem[16'h1ACC] <= 249;
        weight_mem[16'h1ACD] <= 247;
        weight_mem[16'h1ACE] <= 249;
        weight_mem[16'h1ACF] <= 248;
        weight_mem[16'h1AD0] <= 238;
        weight_mem[16'h1AD1] <= 213;
        weight_mem[16'h1AD2] <= 199;
        weight_mem[16'h1AD3] <= 193;
        weight_mem[16'h1AD4] <= 176;
        weight_mem[16'h1AD5] <= 166;
        weight_mem[16'h1AD6] <= 167;
        weight_mem[16'h1AD7] <= 167;
        weight_mem[16'h1AD8] <= 167;
        weight_mem[16'h1AD9] <= 167;
        weight_mem[16'h1ADA] <= 158;
        weight_mem[16'h1ADB] <= 161;
        weight_mem[16'h1ADC] <= 189;
        weight_mem[16'h1ADD] <= 190;
        weight_mem[16'h1ADE] <= 164;
        weight_mem[16'h1ADF] <= 188;
        weight_mem[16'h1AE0] <= 233;
        weight_mem[16'h1AE1] <= 252;
        weight_mem[16'h1AE2] <= 252;
        weight_mem[16'h1AE3] <= 249;
        weight_mem[16'h1AE4] <= 244;
        weight_mem[16'h1AE5] <= 248;
        weight_mem[16'h1AE6] <= 249;
        weight_mem[16'h1AE7] <= 243;
        weight_mem[16'h1AE8] <= 223;
        weight_mem[16'h1AE9] <= 193;
        weight_mem[16'h1AEA] <= 180;
        weight_mem[16'h1AEB] <= 185;
        weight_mem[16'h1AEC] <= 177;
        weight_mem[16'h1AED] <= 167;
        weight_mem[16'h1AEE] <= 167;
        weight_mem[16'h1AEF] <= 167;
        weight_mem[16'h1AF0] <= 167;
        weight_mem[16'h1AF1] <= 167;
        weight_mem[16'h1AF2] <= 158;
        weight_mem[16'h1AF3] <= 158;
        weight_mem[16'h1AF4] <= 183;
        weight_mem[16'h1AF5] <= 148;
        weight_mem[16'h1AF6] <= 158;
        weight_mem[16'h1AF7] <= 198;
        weight_mem[16'h1AF8] <= 225;
        weight_mem[16'h1AF9] <= 243;
        weight_mem[16'h1AFA] <= 252;
        weight_mem[16'h1AFB] <= 252;
        weight_mem[16'h1AFC] <= 251;
        weight_mem[16'h1AFD] <= 252;
        weight_mem[16'h1AFE] <= 253;
        weight_mem[16'h1AFF] <= 245;
        weight_mem[16'h1B00] <= 228;
        weight_mem[16'h1B01] <= 213;
        weight_mem[16'h1B02] <= 199;
        weight_mem[16'h1B03] <= 202;
        weight_mem[16'h1B04] <= 179;
        weight_mem[16'h1B05] <= 167;
        weight_mem[16'h1B06] <= 167;
        weight_mem[16'h1B07] <= 167;
        weight_mem[16'h1B08] <= 167;
        weight_mem[16'h1B09] <= 167;
        weight_mem[16'h1B0A] <= 163;
        weight_mem[16'h1B0B] <= 167;
        weight_mem[16'h1B0C] <= 185;
        weight_mem[16'h1B0D] <= 170;
        weight_mem[16'h1B0E] <= 174;
        weight_mem[16'h1B0F] <= 185;
        weight_mem[16'h1B10] <= 199;
        weight_mem[16'h1B11] <= 217;
        weight_mem[16'h1B12] <= 239;
        weight_mem[16'h1B13] <= 251;
        weight_mem[16'h1B14] <= 253;
        weight_mem[16'h1B15] <= 252;
        weight_mem[16'h1B16] <= 252;
        weight_mem[16'h1B17] <= 243;
        weight_mem[16'h1B18] <= 235;
        weight_mem[16'h1B19] <= 217;
        weight_mem[16'h1B1A] <= 202;
        weight_mem[16'h1B1B] <= 200;
        weight_mem[16'h1B1C] <= 178;
        weight_mem[16'h1B1D] <= 160;
        weight_mem[16'h1B1E] <= 165;
        weight_mem[16'h1B1F] <= 167;
        weight_mem[16'h1B20] <= 167;
        weight_mem[16'h1B21] <= 167;
        weight_mem[16'h1B22] <= 167;
        weight_mem[16'h1B23] <= 180;
        weight_mem[16'h1B24] <= 204;
        weight_mem[16'h1B25] <= 209;
        weight_mem[16'h1B26] <= 190;
        weight_mem[16'h1B27] <= 191;
        weight_mem[16'h1B28] <= 208;
        weight_mem[16'h1B29] <= 229;
        weight_mem[16'h1B2A] <= 235;
        weight_mem[16'h1B2B] <= 245;
        weight_mem[16'h1B2C] <= 249;
        weight_mem[16'h1B2D] <= 245;
        weight_mem[16'h1B2E] <= 242;
        weight_mem[16'h1B2F] <= 244;
        weight_mem[16'h1B30] <= 247;
        weight_mem[16'h1B31] <= 214;
        weight_mem[16'h1B32] <= 197;
        weight_mem[16'h1B33] <= 188;
        weight_mem[16'h1B34] <= 163;
        weight_mem[16'h1B35] <= 145;
        weight_mem[16'h1B36] <= 162;
        weight_mem[16'h1B37] <= 167;
        weight_mem[16'h1B38] <= 167;
        weight_mem[16'h1B39] <= 167;
        weight_mem[16'h1B3A] <= 167;
        weight_mem[16'h1B3B] <= 184;
        weight_mem[16'h1B3C] <= 203;
        weight_mem[16'h1B3D] <= 218;
        weight_mem[16'h1B3E] <= 221;
        weight_mem[16'h1B3F] <= 217;
        weight_mem[16'h1B40] <= 225;
        weight_mem[16'h1B41] <= 236;
        weight_mem[16'h1B42] <= 237;
        weight_mem[16'h1B43] <= 241;
        weight_mem[16'h1B44] <= 242;
        weight_mem[16'h1B45] <= 245;
        weight_mem[16'h1B46] <= 241;
        weight_mem[16'h1B47] <= 241;
        weight_mem[16'h1B48] <= 232;
        weight_mem[16'h1B49] <= 190;
        weight_mem[16'h1B4A] <= 185;
        weight_mem[16'h1B4B] <= 190;
        weight_mem[16'h1B4C] <= 171;
        weight_mem[16'h1B4D] <= 162;
        weight_mem[16'h1B4E] <= 166;
        weight_mem[16'h1B4F] <= 167;
        weight_mem[16'h1B50] <= 167;
        weight_mem[16'h1B51] <= 167;
        weight_mem[16'h1B52] <= 167;
        weight_mem[16'h1B53] <= 173;
        weight_mem[16'h1B54] <= 185;
        weight_mem[16'h1B55] <= 220;
        weight_mem[16'h1B56] <= 238;
        weight_mem[16'h1B57] <= 238;
        weight_mem[16'h1B58] <= 236;
        weight_mem[16'h1B59] <= 238;
        weight_mem[16'h1B5A] <= 241;
        weight_mem[16'h1B5B] <= 245;
        weight_mem[16'h1B5C] <= 248;
        weight_mem[16'h1B5D] <= 245;
        weight_mem[16'h1B5E] <= 237;
        weight_mem[16'h1B5F] <= 230;
        weight_mem[16'h1B60] <= 208;
        weight_mem[16'h1B61] <= 185;
        weight_mem[16'h1B62] <= 192;
        weight_mem[16'h1B63] <= 187;
        weight_mem[16'h1B64] <= 171;
        weight_mem[16'h1B65] <= 167;
        weight_mem[16'h1B66] <= 167;
        weight_mem[16'h1B67] <= 167;
        weight_mem[16'h1B68] <= 167;
        weight_mem[16'h1B69] <= 167;
        weight_mem[16'h1B6A] <= 167;
        weight_mem[16'h1B6B] <= 171;
        weight_mem[16'h1B6C] <= 183;
        weight_mem[16'h1B6D] <= 200;
        weight_mem[16'h1B6E] <= 217;
        weight_mem[16'h1B6F] <= 221;
        weight_mem[16'h1B70] <= 228;
        weight_mem[16'h1B71] <= 228;
        weight_mem[16'h1B72] <= 214;
        weight_mem[16'h1B73] <= 210;
        weight_mem[16'h1B74] <= 227;
        weight_mem[16'h1B75] <= 232;
        weight_mem[16'h1B76] <= 226;
        weight_mem[16'h1B77] <= 217;
        weight_mem[16'h1B78] <= 194;
        weight_mem[16'h1B79] <= 175;
        weight_mem[16'h1B7A] <= 176;
        weight_mem[16'h1B7B] <= 171;
        weight_mem[16'h1B7C] <= 167;
        weight_mem[16'h1B7D] <= 167;
        weight_mem[16'h1B7E] <= 167;
        weight_mem[16'h1B7F] <= 167;
        weight_mem[16'h1B80] <= 167;
        weight_mem[16'h1B81] <= 167;
        weight_mem[16'h1B82] <= 167;
        weight_mem[16'h1B83] <= 173;
        weight_mem[16'h1B84] <= 174;
        weight_mem[16'h1B85] <= 173;
        weight_mem[16'h1B86] <= 176;
        weight_mem[16'h1B87] <= 180;
        weight_mem[16'h1B88] <= 181;
        weight_mem[16'h1B89] <= 179;
        weight_mem[16'h1B8A] <= 166;
        weight_mem[16'h1B8B] <= 162;
        weight_mem[16'h1B8C] <= 161;
        weight_mem[16'h1B8D] <= 194;
        weight_mem[16'h1B8E] <= 192;
        weight_mem[16'h1B8F] <= 182;
        weight_mem[16'h1B90] <= 169;
        weight_mem[16'h1B91] <= 147;
        weight_mem[16'h1B92] <= 161;
        weight_mem[16'h1B93] <= 167;
        weight_mem[16'h1B94] <= 167;
        weight_mem[16'h1B95] <= 167;
        weight_mem[16'h1B96] <= 167;
        weight_mem[16'h1B97] <= 167;
        weight_mem[16'h1B98] <= 167;
        weight_mem[16'h1B99] <= 167;
        weight_mem[16'h1B9A] <= 167;
        weight_mem[16'h1B9B] <= 167;
        weight_mem[16'h1B9C] <= 167;
        weight_mem[16'h1B9D] <= 167;
        weight_mem[16'h1B9E] <= 167;
        weight_mem[16'h1B9F] <= 166;
        weight_mem[16'h1BA0] <= 166;
        weight_mem[16'h1BA1] <= 167;
        weight_mem[16'h1BA2] <= 163;
        weight_mem[16'h1BA3] <= 159;
        weight_mem[16'h1BA4] <= 159;
        weight_mem[16'h1BA5] <= 168;
        weight_mem[16'h1BA6] <= 167;
        weight_mem[16'h1BA7] <= 167;
        weight_mem[16'h1BA8] <= 168;
        weight_mem[16'h1BA9] <= 151;
        weight_mem[16'h1BAA] <= 157;
        weight_mem[16'h1BAB] <= 167;
        weight_mem[16'h1BAC] <= 167;
        weight_mem[16'h1BAD] <= 167;
        weight_mem[16'h1BAE] <= 167;
        weight_mem[16'h1BAF] <= 167;

        // layer 1 neuron 14
        weight_mem[16'h1C00] <= 145;
        weight_mem[16'h1C01] <= 144;
        weight_mem[16'h1C02] <= 145;
        weight_mem[16'h1C03] <= 145;
        weight_mem[16'h1C04] <= 143;
        weight_mem[16'h1C05] <= 144;
        weight_mem[16'h1C06] <= 143;
        weight_mem[16'h1C07] <= 143;
        weight_mem[16'h1C08] <= 143;
        weight_mem[16'h1C09] <= 144;
        weight_mem[16'h1C0A] <= 144;
        weight_mem[16'h1C0B] <= 144;
        weight_mem[16'h1C0C] <= 145;
        weight_mem[16'h1C0D] <= 144;
        weight_mem[16'h1C0E] <= 144;
        weight_mem[16'h1C0F] <= 144;
        weight_mem[16'h1C10] <= 143;
        weight_mem[16'h1C11] <= 144;
        weight_mem[16'h1C12] <= 145;
        weight_mem[16'h1C13] <= 144;
        weight_mem[16'h1C14] <= 143;
        weight_mem[16'h1C15] <= 144;
        weight_mem[16'h1C16] <= 144;
        weight_mem[16'h1C17] <= 143;
        weight_mem[16'h1C18] <= 145;
        weight_mem[16'h1C19] <= 143;
        weight_mem[16'h1C1A] <= 144;
        weight_mem[16'h1C1B] <= 145;
        weight_mem[16'h1C1C] <= 144;
        weight_mem[16'h1C1D] <= 144;
        weight_mem[16'h1C1E] <= 143;
        weight_mem[16'h1C1F] <= 145;
        weight_mem[16'h1C20] <= 145;
        weight_mem[16'h1C21] <= 145;
        weight_mem[16'h1C22] <= 145;
        weight_mem[16'h1C23] <= 147;
        weight_mem[16'h1C24] <= 149;
        weight_mem[16'h1C25] <= 149;
        weight_mem[16'h1C26] <= 145;
        weight_mem[16'h1C27] <= 148;
        weight_mem[16'h1C28] <= 147;
        weight_mem[16'h1C29] <= 149;
        weight_mem[16'h1C2A] <= 148;
        weight_mem[16'h1C2B] <= 144;
        weight_mem[16'h1C2C] <= 143;
        weight_mem[16'h1C2D] <= 142;
        weight_mem[16'h1C2E] <= 145;
        weight_mem[16'h1C2F] <= 144;
        weight_mem[16'h1C30] <= 145;
        weight_mem[16'h1C31] <= 144;
        weight_mem[16'h1C32] <= 145;
        weight_mem[16'h1C33] <= 143;
        weight_mem[16'h1C34] <= 145;
        weight_mem[16'h1C35] <= 145;
        weight_mem[16'h1C36] <= 148;
        weight_mem[16'h1C37] <= 152;
        weight_mem[16'h1C38] <= 153;
        weight_mem[16'h1C39] <= 154;
        weight_mem[16'h1C3A] <= 158;
        weight_mem[16'h1C3B] <= 174;
        weight_mem[16'h1C3C] <= 174;
        weight_mem[16'h1C3D] <= 161;
        weight_mem[16'h1C3E] <= 151;
        weight_mem[16'h1C3F] <= 154;
        weight_mem[16'h1C40] <= 158;
        weight_mem[16'h1C41] <= 156;
        weight_mem[16'h1C42] <= 143;
        weight_mem[16'h1C43] <= 128;
        weight_mem[16'h1C44] <= 134;
        weight_mem[16'h1C45] <= 142;
        weight_mem[16'h1C46] <= 143;
        weight_mem[16'h1C47] <= 143;
        weight_mem[16'h1C48] <= 143;
        weight_mem[16'h1C49] <= 143;
        weight_mem[16'h1C4A] <= 143;
        weight_mem[16'h1C4B] <= 145;
        weight_mem[16'h1C4C] <= 148;
        weight_mem[16'h1C4D] <= 153;
        weight_mem[16'h1C4E] <= 160;
        weight_mem[16'h1C4F] <= 165;
        weight_mem[16'h1C50] <= 166;
        weight_mem[16'h1C51] <= 164;
        weight_mem[16'h1C52] <= 173;
        weight_mem[16'h1C53] <= 197;
        weight_mem[16'h1C54] <= 196;
        weight_mem[16'h1C55] <= 179;
        weight_mem[16'h1C56] <= 176;
        weight_mem[16'h1C57] <= 170;
        weight_mem[16'h1C58] <= 174;
        weight_mem[16'h1C59] <= 165;
        weight_mem[16'h1C5A] <= 148;
        weight_mem[16'h1C5B] <= 131;
        weight_mem[16'h1C5C] <= 139;
        weight_mem[16'h1C5D] <= 145;
        weight_mem[16'h1C5E] <= 146;
        weight_mem[16'h1C5F] <= 144;
        weight_mem[16'h1C60] <= 144;
        weight_mem[16'h1C61] <= 144;
        weight_mem[16'h1C62] <= 143;
        weight_mem[16'h1C63] <= 145;
        weight_mem[16'h1C64] <= 144;
        weight_mem[16'h1C65] <= 151;
        weight_mem[16'h1C66] <= 159;
        weight_mem[16'h1C67] <= 174;
        weight_mem[16'h1C68] <= 191;
        weight_mem[16'h1C69] <= 197;
        weight_mem[16'h1C6A] <= 211;
        weight_mem[16'h1C6B] <= 233;
        weight_mem[16'h1C6C] <= 239;
        weight_mem[16'h1C6D] <= 216;
        weight_mem[16'h1C6E] <= 201;
        weight_mem[16'h1C6F] <= 196;
        weight_mem[16'h1C70] <= 209;
        weight_mem[16'h1C71] <= 219;
        weight_mem[16'h1C72] <= 206;
        weight_mem[16'h1C73] <= 175;
        weight_mem[16'h1C74] <= 156;
        weight_mem[16'h1C75] <= 150;
        weight_mem[16'h1C76] <= 150;
        weight_mem[16'h1C77] <= 144;
        weight_mem[16'h1C78] <= 144;
        weight_mem[16'h1C79] <= 145;
        weight_mem[16'h1C7A] <= 144;
        weight_mem[16'h1C7B] <= 144;
        weight_mem[16'h1C7C] <= 143;
        weight_mem[16'h1C7D] <= 150;
        weight_mem[16'h1C7E] <= 176;
        weight_mem[16'h1C7F] <= 206;
        weight_mem[16'h1C80] <= 231;
        weight_mem[16'h1C81] <= 239;
        weight_mem[16'h1C82] <= 251;
        weight_mem[16'h1C83] <= 254;
        weight_mem[16'h1C84] <= 252;
        weight_mem[16'h1C85] <= 248;
        weight_mem[16'h1C86] <= 246;
        weight_mem[16'h1C87] <= 246;
        weight_mem[16'h1C88] <= 246;
        weight_mem[16'h1C89] <= 235;
        weight_mem[16'h1C8A] <= 207;
        weight_mem[16'h1C8B] <= 175;
        weight_mem[16'h1C8C] <= 142;
        weight_mem[16'h1C8D] <= 144;
        weight_mem[16'h1C8E] <= 145;
        weight_mem[16'h1C8F] <= 144;
        weight_mem[16'h1C90] <= 144;
        weight_mem[16'h1C91] <= 142;
        weight_mem[16'h1C92] <= 142;
        weight_mem[16'h1C93] <= 142;
        weight_mem[16'h1C94] <= 137;
        weight_mem[16'h1C95] <= 150;
        weight_mem[16'h1C96] <= 174;
        weight_mem[16'h1C97] <= 202;
        weight_mem[16'h1C98] <= 234;
        weight_mem[16'h1C99] <= 242;
        weight_mem[16'h1C9A] <= 244;
        weight_mem[16'h1C9B] <= 237;
        weight_mem[16'h1C9C] <= 233;
        weight_mem[16'h1C9D] <= 225;
        weight_mem[16'h1C9E] <= 241;
        weight_mem[16'h1C9F] <= 253;
        weight_mem[16'h1CA0] <= 254;
        weight_mem[16'h1CA1] <= 240;
        weight_mem[16'h1CA2] <= 194;
        weight_mem[16'h1CA3] <= 141;
        weight_mem[16'h1CA4] <= 141;
        weight_mem[16'h1CA5] <= 143;
        weight_mem[16'h1CA6] <= 144;
        weight_mem[16'h1CA7] <= 144;
        weight_mem[16'h1CA8] <= 143;
        weight_mem[16'h1CA9] <= 143;
        weight_mem[16'h1CAA] <= 142;
        weight_mem[16'h1CAB] <= 143;
        weight_mem[16'h1CAC] <= 137;
        weight_mem[16'h1CAD] <= 137;
        weight_mem[16'h1CAE] <= 151;
        weight_mem[16'h1CAF] <= 193;
        weight_mem[16'h1CB0] <= 214;
        weight_mem[16'h1CB1] <= 229;
        weight_mem[16'h1CB2] <= 210;
        weight_mem[16'h1CB3] <= 215;
        weight_mem[16'h1CB4] <= 224;
        weight_mem[16'h1CB5] <= 240;
        weight_mem[16'h1CB6] <= 250;
        weight_mem[16'h1CB7] <= 254;
        weight_mem[16'h1CB8] <= 250;
        weight_mem[16'h1CB9] <= 222;
        weight_mem[16'h1CBA] <= 179;
        weight_mem[16'h1CBB] <= 158;
        weight_mem[16'h1CBC] <= 144;
        weight_mem[16'h1CBD] <= 145;
        weight_mem[16'h1CBE] <= 144;
        weight_mem[16'h1CBF] <= 143;
        weight_mem[16'h1CC0] <= 144;
        weight_mem[16'h1CC1] <= 144;
        weight_mem[16'h1CC2] <= 144;
        weight_mem[16'h1CC3] <= 142;
        weight_mem[16'h1CC4] <= 143;
        weight_mem[16'h1CC5] <= 154;
        weight_mem[16'h1CC6] <= 168;
        weight_mem[16'h1CC7] <= 208;
        weight_mem[16'h1CC8] <= 231;
        weight_mem[16'h1CC9] <= 230;
        weight_mem[16'h1CCA] <= 216;
        weight_mem[16'h1CCB] <= 224;
        weight_mem[16'h1CCC] <= 228;
        weight_mem[16'h1CCD] <= 247;
        weight_mem[16'h1CCE] <= 250;
        weight_mem[16'h1CCF] <= 248;
        weight_mem[16'h1CD0] <= 241;
        weight_mem[16'h1CD1] <= 192;
        weight_mem[16'h1CD2] <= 190;
        weight_mem[16'h1CD3] <= 179;
        weight_mem[16'h1CD4] <= 158;
        weight_mem[16'h1CD5] <= 148;
        weight_mem[16'h1CD6] <= 144;
        weight_mem[16'h1CD7] <= 143;
        weight_mem[16'h1CD8] <= 145;
        weight_mem[16'h1CD9] <= 143;
        weight_mem[16'h1CDA] <= 144;
        weight_mem[16'h1CDB] <= 152;
        weight_mem[16'h1CDC] <= 180;
        weight_mem[16'h1CDD] <= 172;
        weight_mem[16'h1CDE] <= 172;
        weight_mem[16'h1CDF] <= 212;
        weight_mem[16'h1CE0] <= 241;
        weight_mem[16'h1CE1] <= 241;
        weight_mem[16'h1CE2] <= 240;
        weight_mem[16'h1CE3] <= 247;
        weight_mem[16'h1CE4] <= 254;
        weight_mem[16'h1CE5] <= 0;
        weight_mem[16'h1CE6] <= 253;
        weight_mem[16'h1CE7] <= 237;
        weight_mem[16'h1CE8] <= 235;
        weight_mem[16'h1CE9] <= 229;
        weight_mem[16'h1CEA] <= 196;
        weight_mem[16'h1CEB] <= 174;
        weight_mem[16'h1CEC] <= 161;
        weight_mem[16'h1CED] <= 147;
        weight_mem[16'h1CEE] <= 143;
        weight_mem[16'h1CEF] <= 144;
        weight_mem[16'h1CF0] <= 143;
        weight_mem[16'h1CF1] <= 145;
        weight_mem[16'h1CF2] <= 142;
        weight_mem[16'h1CF3] <= 166;
        weight_mem[16'h1CF4] <= 206;
        weight_mem[16'h1CF5] <= 183;
        weight_mem[16'h1CF6] <= 181;
        weight_mem[16'h1CF7] <= 210;
        weight_mem[16'h1CF8] <= 242;
        weight_mem[16'h1CF9] <= 246;
        weight_mem[16'h1CFA] <= 246;
        weight_mem[16'h1CFB] <= 250;
        weight_mem[16'h1CFC] <= 255;
        weight_mem[16'h1CFD] <= 255;
        weight_mem[16'h1CFE] <= 249;
        weight_mem[16'h1CFF] <= 235;
        weight_mem[16'h1D00] <= 242;
        weight_mem[16'h1D01] <= 241;
        weight_mem[16'h1D02] <= 199;
        weight_mem[16'h1D03] <= 168;
        weight_mem[16'h1D04] <= 160;
        weight_mem[16'h1D05] <= 152;
        weight_mem[16'h1D06] <= 145;
        weight_mem[16'h1D07] <= 144;
        weight_mem[16'h1D08] <= 145;
        weight_mem[16'h1D09] <= 143;
        weight_mem[16'h1D0A] <= 144;
        weight_mem[16'h1D0B] <= 164;
        weight_mem[16'h1D0C] <= 206;
        weight_mem[16'h1D0D] <= 224;
        weight_mem[16'h1D0E] <= 231;
        weight_mem[16'h1D0F] <= 235;
        weight_mem[16'h1D10] <= 247;
        weight_mem[16'h1D11] <= 245;
        weight_mem[16'h1D12] <= 240;
        weight_mem[16'h1D13] <= 242;
        weight_mem[16'h1D14] <= 252;
        weight_mem[16'h1D15] <= 249;
        weight_mem[16'h1D16] <= 223;
        weight_mem[16'h1D17] <= 206;
        weight_mem[16'h1D18] <= 219;
        weight_mem[16'h1D19] <= 216;
        weight_mem[16'h1D1A] <= 199;
        weight_mem[16'h1D1B] <= 193;
        weight_mem[16'h1D1C] <= 179;
        weight_mem[16'h1D1D] <= 154;
        weight_mem[16'h1D1E] <= 145;
        weight_mem[16'h1D1F] <= 143;
        weight_mem[16'h1D20] <= 144;
        weight_mem[16'h1D21] <= 143;
        weight_mem[16'h1D22] <= 143;
        weight_mem[16'h1D23] <= 162;
        weight_mem[16'h1D24] <= 188;
        weight_mem[16'h1D25] <= 200;
        weight_mem[16'h1D26] <= 205;
        weight_mem[16'h1D27] <= 211;
        weight_mem[16'h1D28] <= 230;
        weight_mem[16'h1D29] <= 227;
        weight_mem[16'h1D2A] <= 222;
        weight_mem[16'h1D2B] <= 239;
        weight_mem[16'h1D2C] <= 251;
        weight_mem[16'h1D2D] <= 244;
        weight_mem[16'h1D2E] <= 206;
        weight_mem[16'h1D2F] <= 171;
        weight_mem[16'h1D30] <= 180;
        weight_mem[16'h1D31] <= 166;
        weight_mem[16'h1D32] <= 175;
        weight_mem[16'h1D33] <= 193;
        weight_mem[16'h1D34] <= 174;
        weight_mem[16'h1D35] <= 145;
        weight_mem[16'h1D36] <= 144;
        weight_mem[16'h1D37] <= 145;
        weight_mem[16'h1D38] <= 143;
        weight_mem[16'h1D39] <= 144;
        weight_mem[16'h1D3A] <= 144;
        weight_mem[16'h1D3B] <= 150;
        weight_mem[16'h1D3C] <= 158;
        weight_mem[16'h1D3D] <= 157;
        weight_mem[16'h1D3E] <= 179;
        weight_mem[16'h1D3F] <= 203;
        weight_mem[16'h1D40] <= 224;
        weight_mem[16'h1D41] <= 235;
        weight_mem[16'h1D42] <= 225;
        weight_mem[16'h1D43] <= 218;
        weight_mem[16'h1D44] <= 236;
        weight_mem[16'h1D45] <= 236;
        weight_mem[16'h1D46] <= 209;
        weight_mem[16'h1D47] <= 176;
        weight_mem[16'h1D48] <= 154;
        weight_mem[16'h1D49] <= 156;
        weight_mem[16'h1D4A] <= 168;
        weight_mem[16'h1D4B] <= 167;
        weight_mem[16'h1D4C] <= 152;
        weight_mem[16'h1D4D] <= 144;
        weight_mem[16'h1D4E] <= 144;
        weight_mem[16'h1D4F] <= 143;
        weight_mem[16'h1D50] <= 145;
        weight_mem[16'h1D51] <= 144;
        weight_mem[16'h1D52] <= 143;
        weight_mem[16'h1D53] <= 145;
        weight_mem[16'h1D54] <= 139;
        weight_mem[16'h1D55] <= 135;
        weight_mem[16'h1D56] <= 154;
        weight_mem[16'h1D57] <= 184;
        weight_mem[16'h1D58] <= 215;
        weight_mem[16'h1D59] <= 230;
        weight_mem[16'h1D5A] <= 226;
        weight_mem[16'h1D5B] <= 228;
        weight_mem[16'h1D5C] <= 235;
        weight_mem[16'h1D5D] <= 229;
        weight_mem[16'h1D5E] <= 198;
        weight_mem[16'h1D5F] <= 157;
        weight_mem[16'h1D60] <= 150;
        weight_mem[16'h1D61] <= 163;
        weight_mem[16'h1D62] <= 163;
        weight_mem[16'h1D63] <= 162;
        weight_mem[16'h1D64] <= 154;
        weight_mem[16'h1D65] <= 145;
        weight_mem[16'h1D66] <= 144;
        weight_mem[16'h1D67] <= 144;
        weight_mem[16'h1D68] <= 144;
        weight_mem[16'h1D69] <= 144;
        weight_mem[16'h1D6A] <= 144;
        weight_mem[16'h1D6B] <= 145;
        weight_mem[16'h1D6C] <= 144;
        weight_mem[16'h1D6D] <= 145;
        weight_mem[16'h1D6E] <= 154;
        weight_mem[16'h1D6F] <= 185;
        weight_mem[16'h1D70] <= 195;
        weight_mem[16'h1D71] <= 181;
        weight_mem[16'h1D72] <= 168;
        weight_mem[16'h1D73] <= 199;
        weight_mem[16'h1D74] <= 221;
        weight_mem[16'h1D75] <= 201;
        weight_mem[16'h1D76] <= 158;
        weight_mem[16'h1D77] <= 143;
        weight_mem[16'h1D78] <= 143;
        weight_mem[16'h1D79] <= 151;
        weight_mem[16'h1D7A] <= 145;
        weight_mem[16'h1D7B] <= 147;
        weight_mem[16'h1D7C] <= 147;
        weight_mem[16'h1D7D] <= 144;
        weight_mem[16'h1D7E] <= 143;
        weight_mem[16'h1D7F] <= 144;
        weight_mem[16'h1D80] <= 144;
        weight_mem[16'h1D81] <= 145;
        weight_mem[16'h1D82] <= 143;
        weight_mem[16'h1D83] <= 144;
        weight_mem[16'h1D84] <= 144;
        weight_mem[16'h1D85] <= 143;
        weight_mem[16'h1D86] <= 148;
        weight_mem[16'h1D87] <= 162;
        weight_mem[16'h1D88] <= 167;
        weight_mem[16'h1D89] <= 145;
        weight_mem[16'h1D8A] <= 138;
        weight_mem[16'h1D8B] <= 152;
        weight_mem[16'h1D8C] <= 177;
        weight_mem[16'h1D8D] <= 168;
        weight_mem[16'h1D8E] <= 160;
        weight_mem[16'h1D8F] <= 156;
        weight_mem[16'h1D90] <= 140;
        weight_mem[16'h1D91] <= 142;
        weight_mem[16'h1D92] <= 142;
        weight_mem[16'h1D93] <= 143;
        weight_mem[16'h1D94] <= 143;
        weight_mem[16'h1D95] <= 143;
        weight_mem[16'h1D96] <= 144;
        weight_mem[16'h1D97] <= 145;
        weight_mem[16'h1D98] <= 145;
        weight_mem[16'h1D99] <= 143;
        weight_mem[16'h1D9A] <= 144;
        weight_mem[16'h1D9B] <= 143;
        weight_mem[16'h1D9C] <= 144;
        weight_mem[16'h1D9D] <= 144;
        weight_mem[16'h1D9E] <= 144;
        weight_mem[16'h1D9F] <= 144;
        weight_mem[16'h1DA0] <= 145;
        weight_mem[16'h1DA1] <= 144;
        weight_mem[16'h1DA2] <= 143;
        weight_mem[16'h1DA3] <= 145;
        weight_mem[16'h1DA4] <= 145;
        weight_mem[16'h1DA5] <= 151;
        weight_mem[16'h1DA6] <= 153;
        weight_mem[16'h1DA7] <= 151;
        weight_mem[16'h1DA8] <= 144;
        weight_mem[16'h1DA9] <= 146;
        weight_mem[16'h1DAA] <= 145;
        weight_mem[16'h1DAB] <= 143;
        weight_mem[16'h1DAC] <= 144;
        weight_mem[16'h1DAD] <= 144;
        weight_mem[16'h1DAE] <= 143;
        weight_mem[16'h1DAF] <= 145;

        // layer 1 neuron 15
        weight_mem[16'h1E00] <= 185;
        weight_mem[16'h1E01] <= 185;
        weight_mem[16'h1E02] <= 186;
        weight_mem[16'h1E03] <= 186;
        weight_mem[16'h1E04] <= 186;
        weight_mem[16'h1E05] <= 185;
        weight_mem[16'h1E06] <= 186;
        weight_mem[16'h1E07] <= 185;
        weight_mem[16'h1E08] <= 185;
        weight_mem[16'h1E09] <= 185;
        weight_mem[16'h1E0A] <= 186;
        weight_mem[16'h1E0B] <= 184;
        weight_mem[16'h1E0C] <= 185;
        weight_mem[16'h1E0D] <= 186;
        weight_mem[16'h1E0E] <= 185;
        weight_mem[16'h1E0F] <= 186;
        weight_mem[16'h1E10] <= 186;
        weight_mem[16'h1E11] <= 186;
        weight_mem[16'h1E12] <= 184;
        weight_mem[16'h1E13] <= 186;
        weight_mem[16'h1E14] <= 185;
        weight_mem[16'h1E15] <= 185;
        weight_mem[16'h1E16] <= 185;
        weight_mem[16'h1E17] <= 186;
        weight_mem[16'h1E18] <= 186;
        weight_mem[16'h1E19] <= 185;
        weight_mem[16'h1E1A] <= 186;
        weight_mem[16'h1E1B] <= 186;
        weight_mem[16'h1E1C] <= 186;
        weight_mem[16'h1E1D] <= 186;
        weight_mem[16'h1E1E] <= 186;
        weight_mem[16'h1E1F] <= 186;
        weight_mem[16'h1E20] <= 186;
        weight_mem[16'h1E21] <= 186;
        weight_mem[16'h1E22] <= 185;
        weight_mem[16'h1E23] <= 186;
        weight_mem[16'h1E24] <= 188;
        weight_mem[16'h1E25] <= 192;
        weight_mem[16'h1E26] <= 192;
        weight_mem[16'h1E27] <= 194;
        weight_mem[16'h1E28] <= 198;
        weight_mem[16'h1E29] <= 194;
        weight_mem[16'h1E2A] <= 188;
        weight_mem[16'h1E2B] <= 186;
        weight_mem[16'h1E2C] <= 185;
        weight_mem[16'h1E2D] <= 186;
        weight_mem[16'h1E2E] <= 186;
        weight_mem[16'h1E2F] <= 186;
        weight_mem[16'h1E30] <= 186;
        weight_mem[16'h1E31] <= 186;
        weight_mem[16'h1E32] <= 186;
        weight_mem[16'h1E33] <= 186;
        weight_mem[16'h1E34] <= 185;
        weight_mem[16'h1E35] <= 196;
        weight_mem[16'h1E36] <= 200;
        weight_mem[16'h1E37] <= 195;
        weight_mem[16'h1E38] <= 188;
        weight_mem[16'h1E39] <= 192;
        weight_mem[16'h1E3A] <= 196;
        weight_mem[16'h1E3B] <= 211;
        weight_mem[16'h1E3C] <= 223;
        weight_mem[16'h1E3D] <= 223;
        weight_mem[16'h1E3E] <= 220;
        weight_mem[16'h1E3F] <= 215;
        weight_mem[16'h1E40] <= 217;
        weight_mem[16'h1E41] <= 213;
        weight_mem[16'h1E42] <= 191;
        weight_mem[16'h1E43] <= 188;
        weight_mem[16'h1E44] <= 188;
        weight_mem[16'h1E45] <= 186;
        weight_mem[16'h1E46] <= 185;
        weight_mem[16'h1E47] <= 186;
        weight_mem[16'h1E48] <= 185;
        weight_mem[16'h1E49] <= 186;
        weight_mem[16'h1E4A] <= 185;
        weight_mem[16'h1E4B] <= 184;
        weight_mem[16'h1E4C] <= 187;
        weight_mem[16'h1E4D] <= 208;
        weight_mem[16'h1E4E] <= 221;
        weight_mem[16'h1E4F] <= 234;
        weight_mem[16'h1E50] <= 244;
        weight_mem[16'h1E51] <= 249;
        weight_mem[16'h1E52] <= 249;
        weight_mem[16'h1E53] <= 254;
        weight_mem[16'h1E54] <= 255;
        weight_mem[16'h1E55] <= 0;
        weight_mem[16'h1E56] <= 0;
        weight_mem[16'h1E57] <= 253;
        weight_mem[16'h1E58] <= 249;
        weight_mem[16'h1E59] <= 233;
        weight_mem[16'h1E5A] <= 211;
        weight_mem[16'h1E5B] <= 194;
        weight_mem[16'h1E5C] <= 189;
        weight_mem[16'h1E5D] <= 185;
        weight_mem[16'h1E5E] <= 186;
        weight_mem[16'h1E5F] <= 185;
        weight_mem[16'h1E60] <= 186;
        weight_mem[16'h1E61] <= 186;
        weight_mem[16'h1E62] <= 182;
        weight_mem[16'h1E63] <= 179;
        weight_mem[16'h1E64] <= 176;
        weight_mem[16'h1E65] <= 188;
        weight_mem[16'h1E66] <= 224;
        weight_mem[16'h1E67] <= 254;
        weight_mem[16'h1E68] <= 0;
        weight_mem[16'h1E69] <= 254;
        weight_mem[16'h1E6A] <= 0;
        weight_mem[16'h1E6B] <= 2;
        weight_mem[16'h1E6C] <= 1;
        weight_mem[16'h1E6D] <= 1;
        weight_mem[16'h1E6E] <= 1;
        weight_mem[16'h1E6F] <= 0;
        weight_mem[16'h1E70] <= 0;
        weight_mem[16'h1E71] <= 248;
        weight_mem[16'h1E72] <= 221;
        weight_mem[16'h1E73] <= 206;
        weight_mem[16'h1E74] <= 194;
        weight_mem[16'h1E75] <= 186;
        weight_mem[16'h1E76] <= 186;
        weight_mem[16'h1E77] <= 185;
        weight_mem[16'h1E78] <= 185;
        weight_mem[16'h1E79] <= 184;
        weight_mem[16'h1E7A] <= 183;
        weight_mem[16'h1E7B] <= 176;
        weight_mem[16'h1E7C] <= 170;
        weight_mem[16'h1E7D] <= 207;
        weight_mem[16'h1E7E] <= 241;
        weight_mem[16'h1E7F] <= 250;
        weight_mem[16'h1E80] <= 255;
        weight_mem[16'h1E81] <= 1;
        weight_mem[16'h1E82] <= 1;
        weight_mem[16'h1E83] <= 0;
        weight_mem[16'h1E84] <= 0;
        weight_mem[16'h1E85] <= 255;
        weight_mem[16'h1E86] <= 0;
        weight_mem[16'h1E87] <= 0;
        weight_mem[16'h1E88] <= 0;
        weight_mem[16'h1E89] <= 252;
        weight_mem[16'h1E8A] <= 239;
        weight_mem[16'h1E8B] <= 215;
        weight_mem[16'h1E8C] <= 198;
        weight_mem[16'h1E8D] <= 186;
        weight_mem[16'h1E8E] <= 187;
        weight_mem[16'h1E8F] <= 186;
        weight_mem[16'h1E90] <= 185;
        weight_mem[16'h1E91] <= 183;
        weight_mem[16'h1E92] <= 182;
        weight_mem[16'h1E93] <= 184;
        weight_mem[16'h1E94] <= 209;
        weight_mem[16'h1E95] <= 228;
        weight_mem[16'h1E96] <= 226;
        weight_mem[16'h1E97] <= 234;
        weight_mem[16'h1E98] <= 238;
        weight_mem[16'h1E99] <= 253;
        weight_mem[16'h1E9A] <= 255;
        weight_mem[16'h1E9B] <= 254;
        weight_mem[16'h1E9C] <= 252;
        weight_mem[16'h1E9D] <= 252;
        weight_mem[16'h1E9E] <= 0;
        weight_mem[16'h1E9F] <= 0;
        weight_mem[16'h1EA0] <= 0;
        weight_mem[16'h1EA1] <= 251;
        weight_mem[16'h1EA2] <= 229;
        weight_mem[16'h1EA3] <= 208;
        weight_mem[16'h1EA4] <= 203;
        weight_mem[16'h1EA5] <= 190;
        weight_mem[16'h1EA6] <= 185;
        weight_mem[16'h1EA7] <= 185;
        weight_mem[16'h1EA8] <= 184;
        weight_mem[16'h1EA9] <= 182;
        weight_mem[16'h1EAA] <= 184;
        weight_mem[16'h1EAB] <= 185;
        weight_mem[16'h1EAC] <= 220;
        weight_mem[16'h1EAD] <= 230;
        weight_mem[16'h1EAE] <= 216;
        weight_mem[16'h1EAF] <= 228;
        weight_mem[16'h1EB0] <= 229;
        weight_mem[16'h1EB1] <= 249;
        weight_mem[16'h1EB2] <= 254;
        weight_mem[16'h1EB3] <= 250;
        weight_mem[16'h1EB4] <= 237;
        weight_mem[16'h1EB5] <= 251;
        weight_mem[16'h1EB6] <= 0;
        weight_mem[16'h1EB7] <= 0;
        weight_mem[16'h1EB8] <= 3;
        weight_mem[16'h1EB9] <= 252;
        weight_mem[16'h1EBA] <= 230;
        weight_mem[16'h1EBB] <= 191;
        weight_mem[16'h1EBC] <= 193;
        weight_mem[16'h1EBD] <= 193;
        weight_mem[16'h1EBE] <= 185;
        weight_mem[16'h1EBF] <= 185;
        weight_mem[16'h1EC0] <= 185;
        weight_mem[16'h1EC1] <= 185;
        weight_mem[16'h1EC2] <= 188;
        weight_mem[16'h1EC3] <= 184;
        weight_mem[16'h1EC4] <= 208;
        weight_mem[16'h1EC5] <= 246;
        weight_mem[16'h1EC6] <= 241;
        weight_mem[16'h1EC7] <= 241;
        weight_mem[16'h1EC8] <= 254;
        weight_mem[16'h1EC9] <= 0;
        weight_mem[16'h1ECA] <= 0;
        weight_mem[16'h1ECB] <= 243;
        weight_mem[16'h1ECC] <= 254;
        weight_mem[16'h1ECD] <= 0;
        weight_mem[16'h1ECE] <= 0;
        weight_mem[16'h1ECF] <= 0;
        weight_mem[16'h1ED0] <= 0;
        weight_mem[16'h1ED1] <= 246;
        weight_mem[16'h1ED2] <= 216;
        weight_mem[16'h1ED3] <= 175;
        weight_mem[16'h1ED4] <= 183;
        weight_mem[16'h1ED5] <= 186;
        weight_mem[16'h1ED6] <= 185;
        weight_mem[16'h1ED7] <= 184;
        weight_mem[16'h1ED8] <= 185;
        weight_mem[16'h1ED9] <= 184;
        weight_mem[16'h1EDA] <= 192;
        weight_mem[16'h1EDB] <= 199;
        weight_mem[16'h1EDC] <= 187;
        weight_mem[16'h1EDD] <= 202;
        weight_mem[16'h1EDE] <= 223;
        weight_mem[16'h1EDF] <= 241;
        weight_mem[16'h1EE0] <= 250;
        weight_mem[16'h1EE1] <= 0;
        weight_mem[16'h1EE2] <= 0;
        weight_mem[16'h1EE3] <= 254;
        weight_mem[16'h1EE4] <= 0;
        weight_mem[16'h1EE5] <= 0;
        weight_mem[16'h1EE6] <= 0;
        weight_mem[16'h1EE7] <= 254;
        weight_mem[16'h1EE8] <= 250;
        weight_mem[16'h1EE9] <= 248;
        weight_mem[16'h1EEA] <= 202;
        weight_mem[16'h1EEB] <= 174;
        weight_mem[16'h1EEC] <= 188;
        weight_mem[16'h1EED] <= 188;
        weight_mem[16'h1EEE] <= 185;
        weight_mem[16'h1EEF] <= 185;
        weight_mem[16'h1EF0] <= 185;
        weight_mem[16'h1EF1] <= 185;
        weight_mem[16'h1EF2] <= 191;
        weight_mem[16'h1EF3] <= 208;
        weight_mem[16'h1EF4] <= 207;
        weight_mem[16'h1EF5] <= 193;
        weight_mem[16'h1EF6] <= 219;
        weight_mem[16'h1EF7] <= 246;
        weight_mem[16'h1EF8] <= 248;
        weight_mem[16'h1EF9] <= 254;
        weight_mem[16'h1EFA] <= 255;
        weight_mem[16'h1EFB] <= 0;
        weight_mem[16'h1EFC] <= 0;
        weight_mem[16'h1EFD] <= 0;
        weight_mem[16'h1EFE] <= 0;
        weight_mem[16'h1EFF] <= 253;
        weight_mem[16'h1F00] <= 247;
        weight_mem[16'h1F01] <= 244;
        weight_mem[16'h1F02] <= 221;
        weight_mem[16'h1F03] <= 211;
        weight_mem[16'h1F04] <= 200;
        weight_mem[16'h1F05] <= 185;
        weight_mem[16'h1F06] <= 183;
        weight_mem[16'h1F07] <= 184;
        weight_mem[16'h1F08] <= 185;
        weight_mem[16'h1F09] <= 185;
        weight_mem[16'h1F0A] <= 188;
        weight_mem[16'h1F0B] <= 200;
        weight_mem[16'h1F0C] <= 223;
        weight_mem[16'h1F0D] <= 234;
        weight_mem[16'h1F0E] <= 239;
        weight_mem[16'h1F0F] <= 253;
        weight_mem[16'h1F10] <= 254;
        weight_mem[16'h1F11] <= 2;
        weight_mem[16'h1F12] <= 1;
        weight_mem[16'h1F13] <= 255;
        weight_mem[16'h1F14] <= 254;
        weight_mem[16'h1F15] <= 255;
        weight_mem[16'h1F16] <= 253;
        weight_mem[16'h1F17] <= 251;
        weight_mem[16'h1F18] <= 244;
        weight_mem[16'h1F19] <= 245;
        weight_mem[16'h1F1A] <= 229;
        weight_mem[16'h1F1B] <= 222;
        weight_mem[16'h1F1C] <= 221;
        weight_mem[16'h1F1D] <= 195;
        weight_mem[16'h1F1E] <= 181;
        weight_mem[16'h1F1F] <= 184;
        weight_mem[16'h1F20] <= 186;
        weight_mem[16'h1F21] <= 188;
        weight_mem[16'h1F22] <= 190;
        weight_mem[16'h1F23] <= 193;
        weight_mem[16'h1F24] <= 216;
        weight_mem[16'h1F25] <= 239;
        weight_mem[16'h1F26] <= 245;
        weight_mem[16'h1F27] <= 252;
        weight_mem[16'h1F28] <= 254;
        weight_mem[16'h1F29] <= 1;
        weight_mem[16'h1F2A] <= 1;
        weight_mem[16'h1F2B] <= 252;
        weight_mem[16'h1F2C] <= 0;
        weight_mem[16'h1F2D] <= 254;
        weight_mem[16'h1F2E] <= 249;
        weight_mem[16'h1F2F] <= 251;
        weight_mem[16'h1F30] <= 253;
        weight_mem[16'h1F31] <= 248;
        weight_mem[16'h1F32] <= 232;
        weight_mem[16'h1F33] <= 230;
        weight_mem[16'h1F34] <= 226;
        weight_mem[16'h1F35] <= 201;
        weight_mem[16'h1F36] <= 187;
        weight_mem[16'h1F37] <= 186;
        weight_mem[16'h1F38] <= 185;
        weight_mem[16'h1F39] <= 186;
        weight_mem[16'h1F3A] <= 190;
        weight_mem[16'h1F3B] <= 195;
        weight_mem[16'h1F3C] <= 216;
        weight_mem[16'h1F3D] <= 243;
        weight_mem[16'h1F3E] <= 250;
        weight_mem[16'h1F3F] <= 254;
        weight_mem[16'h1F40] <= 0;
        weight_mem[16'h1F41] <= 3;
        weight_mem[16'h1F42] <= 1;
        weight_mem[16'h1F43] <= 255;
        weight_mem[16'h1F44] <= 0;
        weight_mem[16'h1F45] <= 254;
        weight_mem[16'h1F46] <= 254;
        weight_mem[16'h1F47] <= 255;
        weight_mem[16'h1F48] <= 253;
        weight_mem[16'h1F49] <= 253;
        weight_mem[16'h1F4A] <= 245;
        weight_mem[16'h1F4B] <= 228;
        weight_mem[16'h1F4C] <= 202;
        weight_mem[16'h1F4D] <= 190;
        weight_mem[16'h1F4E] <= 186;
        weight_mem[16'h1F4F] <= 186;
        weight_mem[16'h1F50] <= 185;
        weight_mem[16'h1F51] <= 185;
        weight_mem[16'h1F52] <= 186;
        weight_mem[16'h1F53] <= 189;
        weight_mem[16'h1F54] <= 215;
        weight_mem[16'h1F55] <= 237;
        weight_mem[16'h1F56] <= 249;
        weight_mem[16'h1F57] <= 255;
        weight_mem[16'h1F58] <= 2;
        weight_mem[16'h1F59] <= 2;
        weight_mem[16'h1F5A] <= 1;
        weight_mem[16'h1F5B] <= 1;
        weight_mem[16'h1F5C] <= 253;
        weight_mem[16'h1F5D] <= 253;
        weight_mem[16'h1F5E] <= 254;
        weight_mem[16'h1F5F] <= 254;
        weight_mem[16'h1F60] <= 253;
        weight_mem[16'h1F61] <= 253;
        weight_mem[16'h1F62] <= 234;
        weight_mem[16'h1F63] <= 206;
        weight_mem[16'h1F64] <= 185;
        weight_mem[16'h1F65] <= 186;
        weight_mem[16'h1F66] <= 186;
        weight_mem[16'h1F67] <= 186;
        weight_mem[16'h1F68] <= 186;
        weight_mem[16'h1F69] <= 185;
        weight_mem[16'h1F6A] <= 186;
        weight_mem[16'h1F6B] <= 193;
        weight_mem[16'h1F6C] <= 211;
        weight_mem[16'h1F6D] <= 227;
        weight_mem[16'h1F6E] <= 241;
        weight_mem[16'h1F6F] <= 249;
        weight_mem[16'h1F70] <= 0;
        weight_mem[16'h1F71] <= 1;
        weight_mem[16'h1F72] <= 1;
        weight_mem[16'h1F73] <= 250;
        weight_mem[16'h1F74] <= 233;
        weight_mem[16'h1F75] <= 211;
        weight_mem[16'h1F76] <= 234;
        weight_mem[16'h1F77] <= 241;
        weight_mem[16'h1F78] <= 232;
        weight_mem[16'h1F79] <= 217;
        weight_mem[16'h1F7A] <= 208;
        weight_mem[16'h1F7B] <= 203;
        weight_mem[16'h1F7C] <= 187;
        weight_mem[16'h1F7D] <= 185;
        weight_mem[16'h1F7E] <= 185;
        weight_mem[16'h1F7F] <= 185;
        weight_mem[16'h1F80] <= 186;
        weight_mem[16'h1F81] <= 185;
        weight_mem[16'h1F82] <= 186;
        weight_mem[16'h1F83] <= 187;
        weight_mem[16'h1F84] <= 192;
        weight_mem[16'h1F85] <= 204;
        weight_mem[16'h1F86] <= 215;
        weight_mem[16'h1F87] <= 221;
        weight_mem[16'h1F88] <= 235;
        weight_mem[16'h1F89] <= 246;
        weight_mem[16'h1F8A] <= 232;
        weight_mem[16'h1F8B] <= 201;
        weight_mem[16'h1F8C] <= 128;
        weight_mem[16'h1F8D] <= 135;
        weight_mem[16'h1F8E] <= 211;
        weight_mem[16'h1F8F] <= 217;
        weight_mem[16'h1F90] <= 189;
        weight_mem[16'h1F91] <= 182;
        weight_mem[16'h1F92] <= 192;
        weight_mem[16'h1F93] <= 190;
        weight_mem[16'h1F94] <= 185;
        weight_mem[16'h1F95] <= 185;
        weight_mem[16'h1F96] <= 186;
        weight_mem[16'h1F97] <= 186;
        weight_mem[16'h1F98] <= 186;
        weight_mem[16'h1F99] <= 185;
        weight_mem[16'h1F9A] <= 186;
        weight_mem[16'h1F9B] <= 185;
        weight_mem[16'h1F9C] <= 186;
        weight_mem[16'h1F9D] <= 186;
        weight_mem[16'h1F9E] <= 186;
        weight_mem[16'h1F9F] <= 185;
        weight_mem[16'h1FA0] <= 186;
        weight_mem[16'h1FA1] <= 192;
        weight_mem[16'h1FA2] <= 185;
        weight_mem[16'h1FA3] <= 183;
        weight_mem[16'h1FA4] <= 169;
        weight_mem[16'h1FA5] <= 170;
        weight_mem[16'h1FA6] <= 189;
        weight_mem[16'h1FA7] <= 194;
        weight_mem[16'h1FA8] <= 186;
        weight_mem[16'h1FA9] <= 188;
        weight_mem[16'h1FAA] <= 189;
        weight_mem[16'h1FAB] <= 185;
        weight_mem[16'h1FAC] <= 185;
        weight_mem[16'h1FAD] <= 186;
        weight_mem[16'h1FAE] <= 186;
        weight_mem[16'h1FAF] <= 186;

        // layer 1 neuron 16
        weight_mem[16'h2000] <= 1;
        weight_mem[16'h2001] <= 9;
        weight_mem[16'h2002] <= 5;
        weight_mem[16'h2003] <= 2;
        weight_mem[16'h2004] <= 250;
        weight_mem[16'h2005] <= 9;
        weight_mem[16'h2006] <= 254;
        weight_mem[16'h2007] <= 17;
        weight_mem[16'h2008] <= 6;
        weight_mem[16'h2009] <= 7;
        weight_mem[16'h200A] <= 2;
        weight_mem[16'h200B] <= 5;
        weight_mem[16'h200C] <= 251;
        weight_mem[16'h200D] <= 12;
        weight_mem[16'h200E] <= 250;
        weight_mem[16'h200F] <= 5;
        weight_mem[16'h2010] <= 249;
        weight_mem[16'h2011] <= 17;
        weight_mem[16'h2012] <= 12;
        weight_mem[16'h2013] <= 11;
        weight_mem[16'h2014] <= 3;
        weight_mem[16'h2015] <= 1;
        weight_mem[16'h2016] <= 12;
        weight_mem[16'h2017] <= 13;
        weight_mem[16'h2018] <= 255;
        weight_mem[16'h2019] <= 3;
        weight_mem[16'h201A] <= 255;
        weight_mem[16'h201B] <= 14;
        weight_mem[16'h201C] <= 9;
        weight_mem[16'h201D] <= 251;
        weight_mem[16'h201E] <= 13;
        weight_mem[16'h201F] <= 255;
        weight_mem[16'h2020] <= 11;
        weight_mem[16'h2021] <= 254;
        weight_mem[16'h2022] <= 18;
        weight_mem[16'h2023] <= 15;
        weight_mem[16'h2024] <= 11;
        weight_mem[16'h2025] <= 12;
        weight_mem[16'h2026] <= 14;
        weight_mem[16'h2027] <= 14;
        weight_mem[16'h2028] <= 14;
        weight_mem[16'h2029] <= 253;
        weight_mem[16'h202A] <= 19;
        weight_mem[16'h202B] <= 254;
        weight_mem[16'h202C] <= 249;
        weight_mem[16'h202D] <= 252;
        weight_mem[16'h202E] <= 6;
        weight_mem[16'h202F] <= 12;
        weight_mem[16'h2030] <= 9;
        weight_mem[16'h2031] <= 9;
        weight_mem[16'h2032] <= 16;
        weight_mem[16'h2033] <= 6;
        weight_mem[16'h2034] <= 3;
        weight_mem[16'h2035] <= 3;
        weight_mem[16'h2036] <= 253;
        weight_mem[16'h2037] <= 255;
        weight_mem[16'h2038] <= 1;
        weight_mem[16'h2039] <= 11;
        weight_mem[16'h203A] <= 252;
        weight_mem[16'h203B] <= 10;
        weight_mem[16'h203C] <= 3;
        weight_mem[16'h203D] <= 17;
        weight_mem[16'h203E] <= 10;
        weight_mem[16'h203F] <= 8;
        weight_mem[16'h2040] <= 24;
        weight_mem[16'h2041] <= 16;
        weight_mem[16'h2042] <= 2;
        weight_mem[16'h2043] <= 255;
        weight_mem[16'h2044] <= 11;
        weight_mem[16'h2045] <= 2;
        weight_mem[16'h2046] <= 9;
        weight_mem[16'h2047] <= 17;
        weight_mem[16'h2048] <= 252;
        weight_mem[16'h2049] <= 12;
        weight_mem[16'h204A] <= 255;
        weight_mem[16'h204B] <= 255;
        weight_mem[16'h204C] <= 13;
        weight_mem[16'h204D] <= 0;
        weight_mem[16'h204E] <= 3;
        weight_mem[16'h204F] <= 19;
        weight_mem[16'h2050] <= 254;
        weight_mem[16'h2051] <= 233;
        weight_mem[16'h2052] <= 208;
        weight_mem[16'h2053] <= 202;
        weight_mem[16'h2054] <= 220;
        weight_mem[16'h2055] <= 243;
        weight_mem[16'h2056] <= 249;
        weight_mem[16'h2057] <= 255;
        weight_mem[16'h2058] <= 246;
        weight_mem[16'h2059] <= 247;
        weight_mem[16'h205A] <= 0;
        weight_mem[16'h205B] <= 246;
        weight_mem[16'h205C] <= 249;
        weight_mem[16'h205D] <= 0;
        weight_mem[16'h205E] <= 2;
        weight_mem[16'h205F] <= 0;
        weight_mem[16'h2060] <= 17;
        weight_mem[16'h2061] <= 254;
        weight_mem[16'h2062] <= 8;
        weight_mem[16'h2063] <= 10;
        weight_mem[16'h2064] <= 2;
        weight_mem[16'h2065] <= 18;
        weight_mem[16'h2066] <= 2;
        weight_mem[16'h2067] <= 1;
        weight_mem[16'h2068] <= 244;
        weight_mem[16'h2069] <= 229;
        weight_mem[16'h206A] <= 202;
        weight_mem[16'h206B] <= 179;
        weight_mem[16'h206C] <= 193;
        weight_mem[16'h206D] <= 171;
        weight_mem[16'h206E] <= 177;
        weight_mem[16'h206F] <= 197;
        weight_mem[16'h2070] <= 219;
        weight_mem[16'h2071] <= 230;
        weight_mem[16'h2072] <= 246;
        weight_mem[16'h2073] <= 236;
        weight_mem[16'h2074] <= 230;
        weight_mem[16'h2075] <= 243;
        weight_mem[16'h2076] <= 5;
        weight_mem[16'h2077] <= 250;
        weight_mem[16'h2078] <= 249;
        weight_mem[16'h2079] <= 11;
        weight_mem[16'h207A] <= 9;
        weight_mem[16'h207B] <= 10;
        weight_mem[16'h207C] <= 12;
        weight_mem[16'h207D] <= 12;
        weight_mem[16'h207E] <= 10;
        weight_mem[16'h207F] <= 254;
        weight_mem[16'h2080] <= 242;
        weight_mem[16'h2081] <= 233;
        weight_mem[16'h2082] <= 235;
        weight_mem[16'h2083] <= 225;
        weight_mem[16'h2084] <= 1;
        weight_mem[16'h2085] <= 251;
        weight_mem[16'h2086] <= 249;
        weight_mem[16'h2087] <= 233;
        weight_mem[16'h2088] <= 218;
        weight_mem[16'h2089] <= 234;
        weight_mem[16'h208A] <= 233;
        weight_mem[16'h208B] <= 227;
        weight_mem[16'h208C] <= 230;
        weight_mem[16'h208D] <= 225;
        weight_mem[16'h208E] <= 2;
        weight_mem[16'h208F] <= 1;
        weight_mem[16'h2090] <= 16;
        weight_mem[16'h2091] <= 13;
        weight_mem[16'h2092] <= 14;
        weight_mem[16'h2093] <= 25;
        weight_mem[16'h2094] <= 15;
        weight_mem[16'h2095] <= 251;
        weight_mem[16'h2096] <= 242;
        weight_mem[16'h2097] <= 228;
        weight_mem[16'h2098] <= 223;
        weight_mem[16'h2099] <= 238;
        weight_mem[16'h209A] <= 10;
        weight_mem[16'h209B] <= 72;
        weight_mem[16'h209C] <= 78;
        weight_mem[16'h209D] <= 93;
        weight_mem[16'h209E] <= 68;
        weight_mem[16'h209F] <= 37;
        weight_mem[16'h20A0] <= 253;
        weight_mem[16'h20A1] <= 245;
        weight_mem[16'h20A2] <= 245;
        weight_mem[16'h20A3] <= 230;
        weight_mem[16'h20A4] <= 215;
        weight_mem[16'h20A5] <= 223;
        weight_mem[16'h20A6] <= 253;
        weight_mem[16'h20A7] <= 1;
        weight_mem[16'h20A8] <= 249;
        weight_mem[16'h20A9] <= 12;
        weight_mem[16'h20AA] <= 6;
        weight_mem[16'h20AB] <= 20;
        weight_mem[16'h20AC] <= 14;
        weight_mem[16'h20AD] <= 240;
        weight_mem[16'h20AE] <= 230;
        weight_mem[16'h20AF] <= 212;
        weight_mem[16'h20B0] <= 209;
        weight_mem[16'h20B1] <= 227;
        weight_mem[16'h20B2] <= 255;
        weight_mem[16'h20B3] <= 237;
        weight_mem[16'h20B4] <= 204;
        weight_mem[16'h20B5] <= 246;
        weight_mem[16'h20B6] <= 1;
        weight_mem[16'h20B7] <= 2;
        weight_mem[16'h20B8] <= 244;
        weight_mem[16'h20B9] <= 226;
        weight_mem[16'h20BA] <= 209;
        weight_mem[16'h20BB] <= 247;
        weight_mem[16'h20BC] <= 235;
        weight_mem[16'h20BD] <= 253;
        weight_mem[16'h20BE] <= 2;
        weight_mem[16'h20BF] <= 16;
        weight_mem[16'h20C0] <= 17;
        weight_mem[16'h20C1] <= 250;
        weight_mem[16'h20C2] <= 10;
        weight_mem[16'h20C3] <= 5;
        weight_mem[16'h20C4] <= 8;
        weight_mem[16'h20C5] <= 236;
        weight_mem[16'h20C6] <= 235;
        weight_mem[16'h20C7] <= 214;
        weight_mem[16'h20C8] <= 210;
        weight_mem[16'h20C9] <= 231;
        weight_mem[16'h20CA] <= 236;
        weight_mem[16'h20CB] <= 151;
        weight_mem[16'h20CC] <= 128;
        weight_mem[16'h20CD] <= 153;
        weight_mem[16'h20CE] <= 202;
        weight_mem[16'h20CF] <= 230;
        weight_mem[16'h20D0] <= 216;
        weight_mem[16'h20D1] <= 229;
        weight_mem[16'h20D2] <= 252;
        weight_mem[16'h20D3] <= 23;
        weight_mem[16'h20D4] <= 10;
        weight_mem[16'h20D5] <= 250;
        weight_mem[16'h20D6] <= 248;
        weight_mem[16'h20D7] <= 250;
        weight_mem[16'h20D8] <= 13;
        weight_mem[16'h20D9] <= 254;
        weight_mem[16'h20DA] <= 13;
        weight_mem[16'h20DB] <= 6;
        weight_mem[16'h20DC] <= 36;
        weight_mem[16'h20DD] <= 26;
        weight_mem[16'h20DE] <= 15;
        weight_mem[16'h20DF] <= 10;
        weight_mem[16'h20E0] <= 5;
        weight_mem[16'h20E1] <= 237;
        weight_mem[16'h20E2] <= 201;
        weight_mem[16'h20E3] <= 146;
        weight_mem[16'h20E4] <= 153;
        weight_mem[16'h20E5] <= 195;
        weight_mem[16'h20E6] <= 221;
        weight_mem[16'h20E7] <= 234;
        weight_mem[16'h20E8] <= 25;
        weight_mem[16'h20E9] <= 54;
        weight_mem[16'h20EA] <= 52;
        weight_mem[16'h20EB] <= 47;
        weight_mem[16'h20EC] <= 42;
        weight_mem[16'h20ED] <= 17;
        weight_mem[16'h20EE] <= 10;
        weight_mem[16'h20EF] <= 17;
        weight_mem[16'h20F0] <= 8;
        weight_mem[16'h20F1] <= 1;
        weight_mem[16'h20F2] <= 247;
        weight_mem[16'h20F3] <= 16;
        weight_mem[16'h20F4] <= 47;
        weight_mem[16'h20F5] <= 58;
        weight_mem[16'h20F6] <= 55;
        weight_mem[16'h20F7] <= 24;
        weight_mem[16'h20F8] <= 16;
        weight_mem[16'h20F9] <= 255;
        weight_mem[16'h20FA] <= 207;
        weight_mem[16'h20FB] <= 179;
        weight_mem[16'h20FC] <= 210;
        weight_mem[16'h20FD] <= 227;
        weight_mem[16'h20FE] <= 5;
        weight_mem[16'h20FF] <= 58;
        weight_mem[16'h2100] <= 95;
        weight_mem[16'h2101] <= 79;
        weight_mem[16'h2102] <= 48;
        weight_mem[16'h2103] <= 37;
        weight_mem[16'h2104] <= 12;
        weight_mem[16'h2105] <= 22;
        weight_mem[16'h2106] <= 14;
        weight_mem[16'h2107] <= 3;
        weight_mem[16'h2108] <= 6;
        weight_mem[16'h2109] <= 5;
        weight_mem[16'h210A] <= 4;
        weight_mem[16'h210B] <= 24;
        weight_mem[16'h210C] <= 36;
        weight_mem[16'h210D] <= 53;
        weight_mem[16'h210E] <= 48;
        weight_mem[16'h210F] <= 40;
        weight_mem[16'h2110] <= 47;
        weight_mem[16'h2111] <= 51;
        weight_mem[16'h2112] <= 36;
        weight_mem[16'h2113] <= 30;
        weight_mem[16'h2114] <= 27;
        weight_mem[16'h2115] <= 14;
        weight_mem[16'h2116] <= 42;
        weight_mem[16'h2117] <= 65;
        weight_mem[16'h2118] <= 67;
        weight_mem[16'h2119] <= 42;
        weight_mem[16'h211A] <= 41;
        weight_mem[16'h211B] <= 23;
        weight_mem[16'h211C] <= 15;
        weight_mem[16'h211D] <= 19;
        weight_mem[16'h211E] <= 23;
        weight_mem[16'h211F] <= 8;
        weight_mem[16'h2120] <= 16;
        weight_mem[16'h2121] <= 3;
        weight_mem[16'h2122] <= 254;
        weight_mem[16'h2123] <= 254;
        weight_mem[16'h2124] <= 20;
        weight_mem[16'h2125] <= 248;
        weight_mem[16'h2126] <= 18;
        weight_mem[16'h2127] <= 47;
        weight_mem[16'h2128] <= 51;
        weight_mem[16'h2129] <= 90;
        weight_mem[16'h212A] <= 101;
        weight_mem[16'h212B] <= 72;
        weight_mem[16'h212C] <= 35;
        weight_mem[16'h212D] <= 23;
        weight_mem[16'h212E] <= 53;
        weight_mem[16'h212F] <= 44;
        weight_mem[16'h2130] <= 27;
        weight_mem[16'h2131] <= 7;
        weight_mem[16'h2132] <= 12;
        weight_mem[16'h2133] <= 14;
        weight_mem[16'h2134] <= 14;
        weight_mem[16'h2135] <= 15;
        weight_mem[16'h2136] <= 15;
        weight_mem[16'h2137] <= 9;
        weight_mem[16'h2138] <= 254;
        weight_mem[16'h2139] <= 11;
        weight_mem[16'h213A] <= 251;
        weight_mem[16'h213B] <= 11;
        weight_mem[16'h213C] <= 3;
        weight_mem[16'h213D] <= 230;
        weight_mem[16'h213E] <= 217;
        weight_mem[16'h213F] <= 239;
        weight_mem[16'h2140] <= 11;
        weight_mem[16'h2141] <= 41;
        weight_mem[16'h2142] <= 32;
        weight_mem[16'h2143] <= 27;
        weight_mem[16'h2144] <= 15;
        weight_mem[16'h2145] <= 16;
        weight_mem[16'h2146] <= 14;
        weight_mem[16'h2147] <= 19;
        weight_mem[16'h2148] <= 4;
        weight_mem[16'h2149] <= 12;
        weight_mem[16'h214A] <= 8;
        weight_mem[16'h214B] <= 12;
        weight_mem[16'h214C] <= 21;
        weight_mem[16'h214D] <= 19;
        weight_mem[16'h214E] <= 8;
        weight_mem[16'h214F] <= 15;
        weight_mem[16'h2150] <= 254;
        weight_mem[16'h2151] <= 5;
        weight_mem[16'h2152] <= 9;
        weight_mem[16'h2153] <= 253;
        weight_mem[16'h2154] <= 0;
        weight_mem[16'h2155] <= 248;
        weight_mem[16'h2156] <= 227;
        weight_mem[16'h2157] <= 226;
        weight_mem[16'h2158] <= 218;
        weight_mem[16'h2159] <= 206;
        weight_mem[16'h215A] <= 182;
        weight_mem[16'h215B] <= 165;
        weight_mem[16'h215C] <= 177;
        weight_mem[16'h215D] <= 230;
        weight_mem[16'h215E] <= 239;
        weight_mem[16'h215F] <= 253;
        weight_mem[16'h2160] <= 252;
        weight_mem[16'h2161] <= 20;
        weight_mem[16'h2162] <= 23;
        weight_mem[16'h2163] <= 19;
        weight_mem[16'h2164] <= 16;
        weight_mem[16'h2165] <= 16;
        weight_mem[16'h2166] <= 253;
        weight_mem[16'h2167] <= 15;
        weight_mem[16'h2168] <= 12;
        weight_mem[16'h2169] <= 248;
        weight_mem[16'h216A] <= 252;
        weight_mem[16'h216B] <= 250;
        weight_mem[16'h216C] <= 13;
        weight_mem[16'h216D] <= 252;
        weight_mem[16'h216E] <= 5;
        weight_mem[16'h216F] <= 227;
        weight_mem[16'h2170] <= 209;
        weight_mem[16'h2171] <= 186;
        weight_mem[16'h2172] <= 185;
        weight_mem[16'h2173] <= 179;
        weight_mem[16'h2174] <= 194;
        weight_mem[16'h2175] <= 220;
        weight_mem[16'h2176] <= 229;
        weight_mem[16'h2177] <= 232;
        weight_mem[16'h2178] <= 248;
        weight_mem[16'h2179] <= 242;
        weight_mem[16'h217A] <= 4;
        weight_mem[16'h217B] <= 17;
        weight_mem[16'h217C] <= 14;
        weight_mem[16'h217D] <= 18;
        weight_mem[16'h217E] <= 16;
        weight_mem[16'h217F] <= 16;
        weight_mem[16'h2180] <= 253;
        weight_mem[16'h2181] <= 249;
        weight_mem[16'h2182] <= 8;
        weight_mem[16'h2183] <= 10;
        weight_mem[16'h2184] <= 252;
        weight_mem[16'h2185] <= 4;
        weight_mem[16'h2186] <= 246;
        weight_mem[16'h2187] <= 247;
        weight_mem[16'h2188] <= 242;
        weight_mem[16'h2189] <= 242;
        weight_mem[16'h218A] <= 224;
        weight_mem[16'h218B] <= 249;
        weight_mem[16'h218C] <= 236;
        weight_mem[16'h218D] <= 255;
        weight_mem[16'h218E] <= 241;
        weight_mem[16'h218F] <= 231;
        weight_mem[16'h2190] <= 236;
        weight_mem[16'h2191] <= 4;
        weight_mem[16'h2192] <= 245;
        weight_mem[16'h2193] <= 10;
        weight_mem[16'h2194] <= 5;
        weight_mem[16'h2195] <= 10;
        weight_mem[16'h2196] <= 1;
        weight_mem[16'h2197] <= 6;
        weight_mem[16'h2198] <= 13;
        weight_mem[16'h2199] <= 15;
        weight_mem[16'h219A] <= 249;
        weight_mem[16'h219B] <= 254;
        weight_mem[16'h219C] <= 12;
        weight_mem[16'h219D] <= 6;
        weight_mem[16'h219E] <= 6;
        weight_mem[16'h219F] <= 249;
        weight_mem[16'h21A0] <= 4;
        weight_mem[16'h21A1] <= 13;
        weight_mem[16'h21A2] <= 8;
        weight_mem[16'h21A3] <= 255;
        weight_mem[16'h21A4] <= 255;
        weight_mem[16'h21A5] <= 10;
        weight_mem[16'h21A6] <= 250;
        weight_mem[16'h21A7] <= 3;
        weight_mem[16'h21A8] <= 10;
        weight_mem[16'h21A9] <= 255;
        weight_mem[16'h21AA] <= 15;
        weight_mem[16'h21AB] <= 251;
        weight_mem[16'h21AC] <= 11;
        weight_mem[16'h21AD] <= 17;
        weight_mem[16'h21AE] <= 7;
        weight_mem[16'h21AF] <= 9;

        // layer 1 neuron 17
        weight_mem[16'h2200] <= 0;
        weight_mem[16'h2201] <= 0;
        weight_mem[16'h2202] <= 0;
        weight_mem[16'h2203] <= 0;
        weight_mem[16'h2204] <= 0;
        weight_mem[16'h2205] <= 0;
        weight_mem[16'h2206] <= 0;
        weight_mem[16'h2207] <= 0;
        weight_mem[16'h2208] <= 0;
        weight_mem[16'h2209] <= 0;
        weight_mem[16'h220A] <= 0;
        weight_mem[16'h220B] <= 0;
        weight_mem[16'h220C] <= 0;
        weight_mem[16'h220D] <= 0;
        weight_mem[16'h220E] <= 0;
        weight_mem[16'h220F] <= 0;
        weight_mem[16'h2210] <= 0;
        weight_mem[16'h2211] <= 0;
        weight_mem[16'h2212] <= 0;
        weight_mem[16'h2213] <= 0;
        weight_mem[16'h2214] <= 0;
        weight_mem[16'h2215] <= 0;
        weight_mem[16'h2216] <= 0;
        weight_mem[16'h2217] <= 0;
        weight_mem[16'h2218] <= 0;
        weight_mem[16'h2219] <= 0;
        weight_mem[16'h221A] <= 0;
        weight_mem[16'h221B] <= 0;
        weight_mem[16'h221C] <= 0;
        weight_mem[16'h221D] <= 0;
        weight_mem[16'h221E] <= 0;
        weight_mem[16'h221F] <= 0;
        weight_mem[16'h2220] <= 0;
        weight_mem[16'h2221] <= 0;
        weight_mem[16'h2222] <= 0;
        weight_mem[16'h2223] <= 0;
        weight_mem[16'h2224] <= 0;
        weight_mem[16'h2225] <= 0;
        weight_mem[16'h2226] <= 0;
        weight_mem[16'h2227] <= 0;
        weight_mem[16'h2228] <= 0;
        weight_mem[16'h2229] <= 0;
        weight_mem[16'h222A] <= 0;
        weight_mem[16'h222B] <= 0;
        weight_mem[16'h222C] <= 0;
        weight_mem[16'h222D] <= 0;
        weight_mem[16'h222E] <= 0;
        weight_mem[16'h222F] <= 0;
        weight_mem[16'h2230] <= 0;
        weight_mem[16'h2231] <= 0;
        weight_mem[16'h2232] <= 0;
        weight_mem[16'h2233] <= 0;
        weight_mem[16'h2234] <= 0;
        weight_mem[16'h2235] <= 0;
        weight_mem[16'h2236] <= 0;
        weight_mem[16'h2237] <= 0;
        weight_mem[16'h2238] <= 0;
        weight_mem[16'h2239] <= 0;
        weight_mem[16'h223A] <= 0;
        weight_mem[16'h223B] <= 0;
        weight_mem[16'h223C] <= 0;
        weight_mem[16'h223D] <= 0;
        weight_mem[16'h223E] <= 0;
        weight_mem[16'h223F] <= 0;
        weight_mem[16'h2240] <= 0;
        weight_mem[16'h2241] <= 0;
        weight_mem[16'h2242] <= 0;
        weight_mem[16'h2243] <= 0;
        weight_mem[16'h2244] <= 0;
        weight_mem[16'h2245] <= 0;
        weight_mem[16'h2246] <= 0;
        weight_mem[16'h2247] <= 0;
        weight_mem[16'h2248] <= 0;
        weight_mem[16'h2249] <= 0;
        weight_mem[16'h224A] <= 0;
        weight_mem[16'h224B] <= 0;
        weight_mem[16'h224C] <= 0;
        weight_mem[16'h224D] <= 0;
        weight_mem[16'h224E] <= 0;
        weight_mem[16'h224F] <= 0;
        weight_mem[16'h2250] <= 0;
        weight_mem[16'h2251] <= 0;
        weight_mem[16'h2252] <= 0;
        weight_mem[16'h2253] <= 0;
        weight_mem[16'h2254] <= 0;
        weight_mem[16'h2255] <= 0;
        weight_mem[16'h2256] <= 0;
        weight_mem[16'h2257] <= 0;
        weight_mem[16'h2258] <= 0;
        weight_mem[16'h2259] <= 0;
        weight_mem[16'h225A] <= 0;
        weight_mem[16'h225B] <= 0;
        weight_mem[16'h225C] <= 0;
        weight_mem[16'h225D] <= 0;
        weight_mem[16'h225E] <= 0;
        weight_mem[16'h225F] <= 0;
        weight_mem[16'h2260] <= 0;
        weight_mem[16'h2261] <= 0;
        weight_mem[16'h2262] <= 0;
        weight_mem[16'h2263] <= 0;
        weight_mem[16'h2264] <= 0;
        weight_mem[16'h2265] <= 0;
        weight_mem[16'h2266] <= 0;
        weight_mem[16'h2267] <= 0;
        weight_mem[16'h2268] <= 0;
        weight_mem[16'h2269] <= 0;
        weight_mem[16'h226A] <= 0;
        weight_mem[16'h226B] <= 0;
        weight_mem[16'h226C] <= 0;
        weight_mem[16'h226D] <= 0;
        weight_mem[16'h226E] <= 0;
        weight_mem[16'h226F] <= 0;
        weight_mem[16'h2270] <= 0;
        weight_mem[16'h2271] <= 0;
        weight_mem[16'h2272] <= 0;
        weight_mem[16'h2273] <= 0;
        weight_mem[16'h2274] <= 0;
        weight_mem[16'h2275] <= 0;
        weight_mem[16'h2276] <= 0;
        weight_mem[16'h2277] <= 0;
        weight_mem[16'h2278] <= 0;
        weight_mem[16'h2279] <= 0;
        weight_mem[16'h227A] <= 0;
        weight_mem[16'h227B] <= 0;
        weight_mem[16'h227C] <= 0;
        weight_mem[16'h227D] <= 0;
        weight_mem[16'h227E] <= 0;
        weight_mem[16'h227F] <= 0;
        weight_mem[16'h2280] <= 0;
        weight_mem[16'h2281] <= 0;
        weight_mem[16'h2282] <= 0;
        weight_mem[16'h2283] <= 0;
        weight_mem[16'h2284] <= 0;
        weight_mem[16'h2285] <= 0;
        weight_mem[16'h2286] <= 0;
        weight_mem[16'h2287] <= 0;
        weight_mem[16'h2288] <= 0;
        weight_mem[16'h2289] <= 0;
        weight_mem[16'h228A] <= 0;
        weight_mem[16'h228B] <= 0;
        weight_mem[16'h228C] <= 0;
        weight_mem[16'h228D] <= 0;
        weight_mem[16'h228E] <= 0;
        weight_mem[16'h228F] <= 0;
        weight_mem[16'h2290] <= 0;
        weight_mem[16'h2291] <= 0;
        weight_mem[16'h2292] <= 0;
        weight_mem[16'h2293] <= 0;
        weight_mem[16'h2294] <= 0;
        weight_mem[16'h2295] <= 0;
        weight_mem[16'h2296] <= 0;
        weight_mem[16'h2297] <= 0;
        weight_mem[16'h2298] <= 0;
        weight_mem[16'h2299] <= 0;
        weight_mem[16'h229A] <= 0;
        weight_mem[16'h229B] <= 0;
        weight_mem[16'h229C] <= 0;
        weight_mem[16'h229D] <= 0;
        weight_mem[16'h229E] <= 0;
        weight_mem[16'h229F] <= 0;
        weight_mem[16'h22A0] <= 0;
        weight_mem[16'h22A1] <= 0;
        weight_mem[16'h22A2] <= 0;
        weight_mem[16'h22A3] <= 0;
        weight_mem[16'h22A4] <= 0;
        weight_mem[16'h22A5] <= 0;
        weight_mem[16'h22A6] <= 0;
        weight_mem[16'h22A7] <= 0;
        weight_mem[16'h22A8] <= 0;
        weight_mem[16'h22A9] <= 0;
        weight_mem[16'h22AA] <= 0;
        weight_mem[16'h22AB] <= 0;
        weight_mem[16'h22AC] <= 0;
        weight_mem[16'h22AD] <= 0;
        weight_mem[16'h22AE] <= 0;
        weight_mem[16'h22AF] <= 0;
        weight_mem[16'h22B0] <= 0;
        weight_mem[16'h22B1] <= 0;
        weight_mem[16'h22B2] <= 0;
        weight_mem[16'h22B3] <= 0;
        weight_mem[16'h22B4] <= 0;
        weight_mem[16'h22B5] <= 0;
        weight_mem[16'h22B6] <= 0;
        weight_mem[16'h22B7] <= 0;
        weight_mem[16'h22B8] <= 0;
        weight_mem[16'h22B9] <= 0;
        weight_mem[16'h22BA] <= 0;
        weight_mem[16'h22BB] <= 0;
        weight_mem[16'h22BC] <= 0;
        weight_mem[16'h22BD] <= 0;
        weight_mem[16'h22BE] <= 0;
        weight_mem[16'h22BF] <= 0;
        weight_mem[16'h22C0] <= 0;
        weight_mem[16'h22C1] <= 0;
        weight_mem[16'h22C2] <= 0;
        weight_mem[16'h22C3] <= 0;
        weight_mem[16'h22C4] <= 0;
        weight_mem[16'h22C5] <= 0;
        weight_mem[16'h22C6] <= 0;
        weight_mem[16'h22C7] <= 0;
        weight_mem[16'h22C8] <= 0;
        weight_mem[16'h22C9] <= 0;
        weight_mem[16'h22CA] <= 0;
        weight_mem[16'h22CB] <= 0;
        weight_mem[16'h22CC] <= 0;
        weight_mem[16'h22CD] <= 0;
        weight_mem[16'h22CE] <= 0;
        weight_mem[16'h22CF] <= 0;
        weight_mem[16'h22D0] <= 0;
        weight_mem[16'h22D1] <= 0;
        weight_mem[16'h22D2] <= 0;
        weight_mem[16'h22D3] <= 0;
        weight_mem[16'h22D4] <= 0;
        weight_mem[16'h22D5] <= 0;
        weight_mem[16'h22D6] <= 0;
        weight_mem[16'h22D7] <= 0;
        weight_mem[16'h22D8] <= 0;
        weight_mem[16'h22D9] <= 0;
        weight_mem[16'h22DA] <= 0;
        weight_mem[16'h22DB] <= 0;
        weight_mem[16'h22DC] <= 0;
        weight_mem[16'h22DD] <= 0;
        weight_mem[16'h22DE] <= 0;
        weight_mem[16'h22DF] <= 0;
        weight_mem[16'h22E0] <= 0;
        weight_mem[16'h22E1] <= 0;
        weight_mem[16'h22E2] <= 0;
        weight_mem[16'h22E3] <= 0;
        weight_mem[16'h22E4] <= 0;
        weight_mem[16'h22E5] <= 0;
        weight_mem[16'h22E6] <= 0;
        weight_mem[16'h22E7] <= 0;
        weight_mem[16'h22E8] <= 0;
        weight_mem[16'h22E9] <= 0;
        weight_mem[16'h22EA] <= 0;
        weight_mem[16'h22EB] <= 0;
        weight_mem[16'h22EC] <= 0;
        weight_mem[16'h22ED] <= 0;
        weight_mem[16'h22EE] <= 0;
        weight_mem[16'h22EF] <= 0;
        weight_mem[16'h22F0] <= 0;
        weight_mem[16'h22F1] <= 0;
        weight_mem[16'h22F2] <= 0;
        weight_mem[16'h22F3] <= 0;
        weight_mem[16'h22F4] <= 0;
        weight_mem[16'h22F5] <= 0;
        weight_mem[16'h22F6] <= 0;
        weight_mem[16'h22F7] <= 0;
        weight_mem[16'h22F8] <= 0;
        weight_mem[16'h22F9] <= 0;
        weight_mem[16'h22FA] <= 0;
        weight_mem[16'h22FB] <= 0;
        weight_mem[16'h22FC] <= 0;
        weight_mem[16'h22FD] <= 0;
        weight_mem[16'h22FE] <= 0;
        weight_mem[16'h22FF] <= 0;
        weight_mem[16'h2300] <= 0;
        weight_mem[16'h2301] <= 0;
        weight_mem[16'h2302] <= 0;
        weight_mem[16'h2303] <= 0;
        weight_mem[16'h2304] <= 0;
        weight_mem[16'h2305] <= 0;
        weight_mem[16'h2306] <= 0;
        weight_mem[16'h2307] <= 0;
        weight_mem[16'h2308] <= 0;
        weight_mem[16'h2309] <= 0;
        weight_mem[16'h230A] <= 0;
        weight_mem[16'h230B] <= 0;
        weight_mem[16'h230C] <= 0;
        weight_mem[16'h230D] <= 0;
        weight_mem[16'h230E] <= 0;
        weight_mem[16'h230F] <= 0;
        weight_mem[16'h2310] <= 0;
        weight_mem[16'h2311] <= 0;
        weight_mem[16'h2312] <= 0;
        weight_mem[16'h2313] <= 0;
        weight_mem[16'h2314] <= 0;
        weight_mem[16'h2315] <= 0;
        weight_mem[16'h2316] <= 0;
        weight_mem[16'h2317] <= 0;
        weight_mem[16'h2318] <= 0;
        weight_mem[16'h2319] <= 0;
        weight_mem[16'h231A] <= 0;
        weight_mem[16'h231B] <= 0;
        weight_mem[16'h231C] <= 0;
        weight_mem[16'h231D] <= 0;
        weight_mem[16'h231E] <= 0;
        weight_mem[16'h231F] <= 0;
        weight_mem[16'h2320] <= 0;
        weight_mem[16'h2321] <= 0;
        weight_mem[16'h2322] <= 0;
        weight_mem[16'h2323] <= 0;
        weight_mem[16'h2324] <= 0;
        weight_mem[16'h2325] <= 0;
        weight_mem[16'h2326] <= 0;
        weight_mem[16'h2327] <= 0;
        weight_mem[16'h2328] <= 0;
        weight_mem[16'h2329] <= 0;
        weight_mem[16'h232A] <= 0;
        weight_mem[16'h232B] <= 0;
        weight_mem[16'h232C] <= 0;
        weight_mem[16'h232D] <= 0;
        weight_mem[16'h232E] <= 0;
        weight_mem[16'h232F] <= 0;
        weight_mem[16'h2330] <= 0;
        weight_mem[16'h2331] <= 0;
        weight_mem[16'h2332] <= 0;
        weight_mem[16'h2333] <= 0;
        weight_mem[16'h2334] <= 0;
        weight_mem[16'h2335] <= 0;
        weight_mem[16'h2336] <= 0;
        weight_mem[16'h2337] <= 0;
        weight_mem[16'h2338] <= 0;
        weight_mem[16'h2339] <= 0;
        weight_mem[16'h233A] <= 0;
        weight_mem[16'h233B] <= 0;
        weight_mem[16'h233C] <= 0;
        weight_mem[16'h233D] <= 0;
        weight_mem[16'h233E] <= 0;
        weight_mem[16'h233F] <= 0;
        weight_mem[16'h2340] <= 0;
        weight_mem[16'h2341] <= 0;
        weight_mem[16'h2342] <= 0;
        weight_mem[16'h2343] <= 0;
        weight_mem[16'h2344] <= 0;
        weight_mem[16'h2345] <= 0;
        weight_mem[16'h2346] <= 0;
        weight_mem[16'h2347] <= 0;
        weight_mem[16'h2348] <= 0;
        weight_mem[16'h2349] <= 0;
        weight_mem[16'h234A] <= 0;
        weight_mem[16'h234B] <= 0;
        weight_mem[16'h234C] <= 0;
        weight_mem[16'h234D] <= 0;
        weight_mem[16'h234E] <= 0;
        weight_mem[16'h234F] <= 0;
        weight_mem[16'h2350] <= 0;
        weight_mem[16'h2351] <= 0;
        weight_mem[16'h2352] <= 0;
        weight_mem[16'h2353] <= 0;
        weight_mem[16'h2354] <= 0;
        weight_mem[16'h2355] <= 0;
        weight_mem[16'h2356] <= 0;
        weight_mem[16'h2357] <= 0;
        weight_mem[16'h2358] <= 0;
        weight_mem[16'h2359] <= 0;
        weight_mem[16'h235A] <= 0;
        weight_mem[16'h235B] <= 0;
        weight_mem[16'h235C] <= 0;
        weight_mem[16'h235D] <= 0;
        weight_mem[16'h235E] <= 0;
        weight_mem[16'h235F] <= 0;
        weight_mem[16'h2360] <= 0;
        weight_mem[16'h2361] <= 0;
        weight_mem[16'h2362] <= 0;
        weight_mem[16'h2363] <= 0;
        weight_mem[16'h2364] <= 0;
        weight_mem[16'h2365] <= 0;
        weight_mem[16'h2366] <= 0;
        weight_mem[16'h2367] <= 0;
        weight_mem[16'h2368] <= 0;
        weight_mem[16'h2369] <= 0;
        weight_mem[16'h236A] <= 0;
        weight_mem[16'h236B] <= 0;
        weight_mem[16'h236C] <= 0;
        weight_mem[16'h236D] <= 0;
        weight_mem[16'h236E] <= 0;
        weight_mem[16'h236F] <= 0;
        weight_mem[16'h2370] <= 0;
        weight_mem[16'h2371] <= 0;
        weight_mem[16'h2372] <= 0;
        weight_mem[16'h2373] <= 0;
        weight_mem[16'h2374] <= 0;
        weight_mem[16'h2375] <= 0;
        weight_mem[16'h2376] <= 0;
        weight_mem[16'h2377] <= 0;
        weight_mem[16'h2378] <= 0;
        weight_mem[16'h2379] <= 0;
        weight_mem[16'h237A] <= 0;
        weight_mem[16'h237B] <= 0;
        weight_mem[16'h237C] <= 0;
        weight_mem[16'h237D] <= 0;
        weight_mem[16'h237E] <= 0;
        weight_mem[16'h237F] <= 0;
        weight_mem[16'h2380] <= 0;
        weight_mem[16'h2381] <= 0;
        weight_mem[16'h2382] <= 0;
        weight_mem[16'h2383] <= 0;
        weight_mem[16'h2384] <= 0;
        weight_mem[16'h2385] <= 0;
        weight_mem[16'h2386] <= 0;
        weight_mem[16'h2387] <= 0;
        weight_mem[16'h2388] <= 0;
        weight_mem[16'h2389] <= 0;
        weight_mem[16'h238A] <= 0;
        weight_mem[16'h238B] <= 0;
        weight_mem[16'h238C] <= 0;
        weight_mem[16'h238D] <= 0;
        weight_mem[16'h238E] <= 0;
        weight_mem[16'h238F] <= 0;
        weight_mem[16'h2390] <= 0;
        weight_mem[16'h2391] <= 0;
        weight_mem[16'h2392] <= 0;
        weight_mem[16'h2393] <= 0;
        weight_mem[16'h2394] <= 0;
        weight_mem[16'h2395] <= 0;
        weight_mem[16'h2396] <= 0;
        weight_mem[16'h2397] <= 0;
        weight_mem[16'h2398] <= 0;
        weight_mem[16'h2399] <= 0;
        weight_mem[16'h239A] <= 0;
        weight_mem[16'h239B] <= 0;
        weight_mem[16'h239C] <= 0;
        weight_mem[16'h239D] <= 0;
        weight_mem[16'h239E] <= 0;
        weight_mem[16'h239F] <= 0;
        weight_mem[16'h23A0] <= 0;
        weight_mem[16'h23A1] <= 0;
        weight_mem[16'h23A2] <= 0;
        weight_mem[16'h23A3] <= 0;
        weight_mem[16'h23A4] <= 0;
        weight_mem[16'h23A5] <= 0;
        weight_mem[16'h23A6] <= 0;
        weight_mem[16'h23A7] <= 0;
        weight_mem[16'h23A8] <= 0;
        weight_mem[16'h23A9] <= 0;
        weight_mem[16'h23AA] <= 0;
        weight_mem[16'h23AB] <= 0;
        weight_mem[16'h23AC] <= 0;
        weight_mem[16'h23AD] <= 0;
        weight_mem[16'h23AE] <= 0;
        weight_mem[16'h23AF] <= 0;

        // layer 1 neuron 18
        weight_mem[16'h2400] <= 161;
        weight_mem[16'h2401] <= 161;
        weight_mem[16'h2402] <= 161;
        weight_mem[16'h2403] <= 161;
        weight_mem[16'h2404] <= 161;
        weight_mem[16'h2405] <= 161;
        weight_mem[16'h2406] <= 161;
        weight_mem[16'h2407] <= 161;
        weight_mem[16'h2408] <= 161;
        weight_mem[16'h2409] <= 161;
        weight_mem[16'h240A] <= 161;
        weight_mem[16'h240B] <= 161;
        weight_mem[16'h240C] <= 161;
        weight_mem[16'h240D] <= 161;
        weight_mem[16'h240E] <= 161;
        weight_mem[16'h240F] <= 161;
        weight_mem[16'h2410] <= 161;
        weight_mem[16'h2411] <= 161;
        weight_mem[16'h2412] <= 161;
        weight_mem[16'h2413] <= 161;
        weight_mem[16'h2414] <= 161;
        weight_mem[16'h2415] <= 161;
        weight_mem[16'h2416] <= 161;
        weight_mem[16'h2417] <= 161;
        weight_mem[16'h2418] <= 161;
        weight_mem[16'h2419] <= 161;
        weight_mem[16'h241A] <= 161;
        weight_mem[16'h241B] <= 161;
        weight_mem[16'h241C] <= 161;
        weight_mem[16'h241D] <= 161;
        weight_mem[16'h241E] <= 161;
        weight_mem[16'h241F] <= 161;
        weight_mem[16'h2420] <= 161;
        weight_mem[16'h2421] <= 161;
        weight_mem[16'h2422] <= 161;
        weight_mem[16'h2423] <= 161;
        weight_mem[16'h2424] <= 160;
        weight_mem[16'h2425] <= 162;
        weight_mem[16'h2426] <= 162;
        weight_mem[16'h2427] <= 162;
        weight_mem[16'h2428] <= 162;
        weight_mem[16'h2429] <= 162;
        weight_mem[16'h242A] <= 162;
        weight_mem[16'h242B] <= 161;
        weight_mem[16'h242C] <= 161;
        weight_mem[16'h242D] <= 161;
        weight_mem[16'h242E] <= 161;
        weight_mem[16'h242F] <= 161;
        weight_mem[16'h2430] <= 161;
        weight_mem[16'h2431] <= 161;
        weight_mem[16'h2432] <= 161;
        weight_mem[16'h2433] <= 161;
        weight_mem[16'h2434] <= 161;
        weight_mem[16'h2435] <= 161;
        weight_mem[16'h2436] <= 161;
        weight_mem[16'h2437] <= 161;
        weight_mem[16'h2438] <= 161;
        weight_mem[16'h2439] <= 160;
        weight_mem[16'h243A] <= 159;
        weight_mem[16'h243B] <= 157;
        weight_mem[16'h243C] <= 157;
        weight_mem[16'h243D] <= 175;
        weight_mem[16'h243E] <= 173;
        weight_mem[16'h243F] <= 171;
        weight_mem[16'h2440] <= 170;
        weight_mem[16'h2441] <= 171;
        weight_mem[16'h2442] <= 166;
        weight_mem[16'h2443] <= 162;
        weight_mem[16'h2444] <= 161;
        weight_mem[16'h2445] <= 161;
        weight_mem[16'h2446] <= 161;
        weight_mem[16'h2447] <= 161;
        weight_mem[16'h2448] <= 161;
        weight_mem[16'h2449] <= 161;
        weight_mem[16'h244A] <= 161;
        weight_mem[16'h244B] <= 161;
        weight_mem[16'h244C] <= 160;
        weight_mem[16'h244D] <= 160;
        weight_mem[16'h244E] <= 160;
        weight_mem[16'h244F] <= 159;
        weight_mem[16'h2450] <= 154;
        weight_mem[16'h2451] <= 151;
        weight_mem[16'h2452] <= 147;
        weight_mem[16'h2453] <= 136;
        weight_mem[16'h2454] <= 158;
        weight_mem[16'h2455] <= 182;
        weight_mem[16'h2456] <= 180;
        weight_mem[16'h2457] <= 183;
        weight_mem[16'h2458] <= 176;
        weight_mem[16'h2459] <= 182;
        weight_mem[16'h245A] <= 174;
        weight_mem[16'h245B] <= 164;
        weight_mem[16'h245C] <= 162;
        weight_mem[16'h245D] <= 161;
        weight_mem[16'h245E] <= 161;
        weight_mem[16'h245F] <= 161;
        weight_mem[16'h2460] <= 161;
        weight_mem[16'h2461] <= 161;
        weight_mem[16'h2462] <= 161;
        weight_mem[16'h2463] <= 161;
        weight_mem[16'h2464] <= 161;
        weight_mem[16'h2465] <= 162;
        weight_mem[16'h2466] <= 168;
        weight_mem[16'h2467] <= 166;
        weight_mem[16'h2468] <= 153;
        weight_mem[16'h2469] <= 151;
        weight_mem[16'h246A] <= 143;
        weight_mem[16'h246B] <= 128;
        weight_mem[16'h246C] <= 173;
        weight_mem[16'h246D] <= 184;
        weight_mem[16'h246E] <= 171;
        weight_mem[16'h246F] <= 174;
        weight_mem[16'h2470] <= 160;
        weight_mem[16'h2471] <= 158;
        weight_mem[16'h2472] <= 165;
        weight_mem[16'h2473] <= 158;
        weight_mem[16'h2474] <= 163;
        weight_mem[16'h2475] <= 162;
        weight_mem[16'h2476] <= 162;
        weight_mem[16'h2477] <= 161;
        weight_mem[16'h2478] <= 161;
        weight_mem[16'h2479] <= 161;
        weight_mem[16'h247A] <= 161;
        weight_mem[16'h247B] <= 161;
        weight_mem[16'h247C] <= 161;
        weight_mem[16'h247D] <= 169;
        weight_mem[16'h247E] <= 181;
        weight_mem[16'h247F] <= 170;
        weight_mem[16'h2480] <= 163;
        weight_mem[16'h2481] <= 180;
        weight_mem[16'h2482] <= 196;
        weight_mem[16'h2483] <= 210;
        weight_mem[16'h2484] <= 225;
        weight_mem[16'h2485] <= 204;
        weight_mem[16'h2486] <= 193;
        weight_mem[16'h2487] <= 203;
        weight_mem[16'h2488] <= 182;
        weight_mem[16'h2489] <= 158;
        weight_mem[16'h248A] <= 158;
        weight_mem[16'h248B] <= 163;
        weight_mem[16'h248C] <= 166;
        weight_mem[16'h248D] <= 164;
        weight_mem[16'h248E] <= 163;
        weight_mem[16'h248F] <= 161;
        weight_mem[16'h2490] <= 161;
        weight_mem[16'h2491] <= 161;
        weight_mem[16'h2492] <= 162;
        weight_mem[16'h2493] <= 162;
        weight_mem[16'h2494] <= 165;
        weight_mem[16'h2495] <= 171;
        weight_mem[16'h2496] <= 171;
        weight_mem[16'h2497] <= 166;
        weight_mem[16'h2498] <= 158;
        weight_mem[16'h2499] <= 182;
        weight_mem[16'h249A] <= 203;
        weight_mem[16'h249B] <= 219;
        weight_mem[16'h249C] <= 223;
        weight_mem[16'h249D] <= 214;
        weight_mem[16'h249E] <= 223;
        weight_mem[16'h249F] <= 230;
        weight_mem[16'h24A0] <= 200;
        weight_mem[16'h24A1] <= 166;
        weight_mem[16'h24A2] <= 157;
        weight_mem[16'h24A3] <= 166;
        weight_mem[16'h24A4] <= 166;
        weight_mem[16'h24A5] <= 165;
        weight_mem[16'h24A6] <= 163;
        weight_mem[16'h24A7] <= 161;
        weight_mem[16'h24A8] <= 161;
        weight_mem[16'h24A9] <= 161;
        weight_mem[16'h24AA] <= 161;
        weight_mem[16'h24AB] <= 162;
        weight_mem[16'h24AC] <= 167;
        weight_mem[16'h24AD] <= 169;
        weight_mem[16'h24AE] <= 169;
        weight_mem[16'h24AF] <= 171;
        weight_mem[16'h24B0] <= 149;
        weight_mem[16'h24B1] <= 161;
        weight_mem[16'h24B2] <= 166;
        weight_mem[16'h24B3] <= 188;
        weight_mem[16'h24B4] <= 209;
        weight_mem[16'h24B5] <= 219;
        weight_mem[16'h24B6] <= 214;
        weight_mem[16'h24B7] <= 217;
        weight_mem[16'h24B8] <= 199;
        weight_mem[16'h24B9] <= 174;
        weight_mem[16'h24BA] <= 158;
        weight_mem[16'h24BB] <= 162;
        weight_mem[16'h24BC] <= 166;
        weight_mem[16'h24BD] <= 164;
        weight_mem[16'h24BE] <= 162;
        weight_mem[16'h24BF] <= 161;
        weight_mem[16'h24C0] <= 161;
        weight_mem[16'h24C1] <= 161;
        weight_mem[16'h24C2] <= 161;
        weight_mem[16'h24C3] <= 161;
        weight_mem[16'h24C4] <= 163;
        weight_mem[16'h24C5] <= 165;
        weight_mem[16'h24C6] <= 170;
        weight_mem[16'h24C7] <= 183;
        weight_mem[16'h24C8] <= 172;
        weight_mem[16'h24C9] <= 157;
        weight_mem[16'h24CA] <= 156;
        weight_mem[16'h24CB] <= 186;
        weight_mem[16'h24CC] <= 205;
        weight_mem[16'h24CD] <= 194;
        weight_mem[16'h24CE] <= 169;
        weight_mem[16'h24CF] <= 167;
        weight_mem[16'h24D0] <= 183;
        weight_mem[16'h24D1] <= 191;
        weight_mem[16'h24D2] <= 173;
        weight_mem[16'h24D3] <= 159;
        weight_mem[16'h24D4] <= 163;
        weight_mem[16'h24D5] <= 162;
        weight_mem[16'h24D6] <= 161;
        weight_mem[16'h24D7] <= 161;
        weight_mem[16'h24D8] <= 161;
        weight_mem[16'h24D9] <= 161;
        weight_mem[16'h24DA] <= 161;
        weight_mem[16'h24DB] <= 162;
        weight_mem[16'h24DC] <= 161;
        weight_mem[16'h24DD] <= 161;
        weight_mem[16'h24DE] <= 169;
        weight_mem[16'h24DF] <= 189;
        weight_mem[16'h24E0] <= 180;
        weight_mem[16'h24E1] <= 155;
        weight_mem[16'h24E2] <= 164;
        weight_mem[16'h24E3] <= 176;
        weight_mem[16'h24E4] <= 186;
        weight_mem[16'h24E5] <= 192;
        weight_mem[16'h24E6] <= 170;
        weight_mem[16'h24E7] <= 156;
        weight_mem[16'h24E8] <= 161;
        weight_mem[16'h24E9] <= 182;
        weight_mem[16'h24EA] <= 175;
        weight_mem[16'h24EB] <= 157;
        weight_mem[16'h24EC] <= 160;
        weight_mem[16'h24ED] <= 162;
        weight_mem[16'h24EE] <= 161;
        weight_mem[16'h24EF] <= 161;
        weight_mem[16'h24F0] <= 161;
        weight_mem[16'h24F1] <= 161;
        weight_mem[16'h24F2] <= 162;
        weight_mem[16'h24F3] <= 162;
        weight_mem[16'h24F4] <= 164;
        weight_mem[16'h24F5] <= 162;
        weight_mem[16'h24F6] <= 164;
        weight_mem[16'h24F7] <= 176;
        weight_mem[16'h24F8] <= 168;
        weight_mem[16'h24F9] <= 175;
        weight_mem[16'h24FA] <= 175;
        weight_mem[16'h24FB] <= 170;
        weight_mem[16'h24FC] <= 186;
        weight_mem[16'h24FD] <= 187;
        weight_mem[16'h24FE] <= 157;
        weight_mem[16'h24FF] <= 140;
        weight_mem[16'h2500] <= 146;
        weight_mem[16'h2501] <= 172;
        weight_mem[16'h2502] <= 180;
        weight_mem[16'h2503] <= 166;
        weight_mem[16'h2504] <= 161;
        weight_mem[16'h2505] <= 161;
        weight_mem[16'h2506] <= 162;
        weight_mem[16'h2507] <= 161;
        weight_mem[16'h2508] <= 161;
        weight_mem[16'h2509] <= 161;
        weight_mem[16'h250A] <= 162;
        weight_mem[16'h250B] <= 166;
        weight_mem[16'h250C] <= 174;
        weight_mem[16'h250D] <= 170;
        weight_mem[16'h250E] <= 161;
        weight_mem[16'h250F] <= 167;
        weight_mem[16'h2510] <= 177;
        weight_mem[16'h2511] <= 179;
        weight_mem[16'h2512] <= 182;
        weight_mem[16'h2513] <= 169;
        weight_mem[16'h2514] <= 191;
        weight_mem[16'h2515] <= 179;
        weight_mem[16'h2516] <= 142;
        weight_mem[16'h2517] <= 140;
        weight_mem[16'h2518] <= 150;
        weight_mem[16'h2519] <= 180;
        weight_mem[16'h251A] <= 182;
        weight_mem[16'h251B] <= 176;
        weight_mem[16'h251C] <= 165;
        weight_mem[16'h251D] <= 162;
        weight_mem[16'h251E] <= 162;
        weight_mem[16'h251F] <= 162;
        weight_mem[16'h2520] <= 161;
        weight_mem[16'h2521] <= 161;
        weight_mem[16'h2522] <= 162;
        weight_mem[16'h2523] <= 171;
        weight_mem[16'h2524] <= 179;
        weight_mem[16'h2525] <= 178;
        weight_mem[16'h2526] <= 167;
        weight_mem[16'h2527] <= 170;
        weight_mem[16'h2528] <= 175;
        weight_mem[16'h2529] <= 181;
        weight_mem[16'h252A] <= 166;
        weight_mem[16'h252B] <= 167;
        weight_mem[16'h252C] <= 205;
        weight_mem[16'h252D] <= 184;
        weight_mem[16'h252E] <= 145;
        weight_mem[16'h252F] <= 156;
        weight_mem[16'h2530] <= 174;
        weight_mem[16'h2531] <= 176;
        weight_mem[16'h2532] <= 171;
        weight_mem[16'h2533] <= 180;
        weight_mem[16'h2534] <= 169;
        weight_mem[16'h2535] <= 162;
        weight_mem[16'h2536] <= 162;
        weight_mem[16'h2537] <= 162;
        weight_mem[16'h2538] <= 161;
        weight_mem[16'h2539] <= 161;
        weight_mem[16'h253A] <= 161;
        weight_mem[16'h253B] <= 166;
        weight_mem[16'h253C] <= 177;
        weight_mem[16'h253D] <= 179;
        weight_mem[16'h253E] <= 174;
        weight_mem[16'h253F] <= 183;
        weight_mem[16'h2540] <= 172;
        weight_mem[16'h2541] <= 160;
        weight_mem[16'h2542] <= 171;
        weight_mem[16'h2543] <= 173;
        weight_mem[16'h2544] <= 198;
        weight_mem[16'h2545] <= 156;
        weight_mem[16'h2546] <= 143;
        weight_mem[16'h2547] <= 166;
        weight_mem[16'h2548] <= 168;
        weight_mem[16'h2549] <= 157;
        weight_mem[16'h254A] <= 161;
        weight_mem[16'h254B] <= 177;
        weight_mem[16'h254C] <= 167;
        weight_mem[16'h254D] <= 162;
        weight_mem[16'h254E] <= 162;
        weight_mem[16'h254F] <= 161;
        weight_mem[16'h2550] <= 161;
        weight_mem[16'h2551] <= 161;
        weight_mem[16'h2552] <= 161;
        weight_mem[16'h2553] <= 163;
        weight_mem[16'h2554] <= 169;
        weight_mem[16'h2555] <= 170;
        weight_mem[16'h2556] <= 167;
        weight_mem[16'h2557] <= 182;
        weight_mem[16'h2558] <= 176;
        weight_mem[16'h2559] <= 176;
        weight_mem[16'h255A] <= 180;
        weight_mem[16'h255B] <= 175;
        weight_mem[16'h255C] <= 164;
        weight_mem[16'h255D] <= 137;
        weight_mem[16'h255E] <= 151;
        weight_mem[16'h255F] <= 153;
        weight_mem[16'h2560] <= 145;
        weight_mem[16'h2561] <= 148;
        weight_mem[16'h2562] <= 159;
        weight_mem[16'h2563] <= 173;
        weight_mem[16'h2564] <= 168;
        weight_mem[16'h2565] <= 161;
        weight_mem[16'h2566] <= 161;
        weight_mem[16'h2567] <= 161;
        weight_mem[16'h2568] <= 161;
        weight_mem[16'h2569] <= 161;
        weight_mem[16'h256A] <= 161;
        weight_mem[16'h256B] <= 163;
        weight_mem[16'h256C] <= 166;
        weight_mem[16'h256D] <= 165;
        weight_mem[16'h256E] <= 163;
        weight_mem[16'h256F] <= 174;
        weight_mem[16'h2570] <= 176;
        weight_mem[16'h2571] <= 174;
        weight_mem[16'h2572] <= 173;
        weight_mem[16'h2573] <= 173;
        weight_mem[16'h2574] <= 162;
        weight_mem[16'h2575] <= 153;
        weight_mem[16'h2576] <= 159;
        weight_mem[16'h2577] <= 158;
        weight_mem[16'h2578] <= 158;
        weight_mem[16'h2579] <= 161;
        weight_mem[16'h257A] <= 164;
        weight_mem[16'h257B] <= 173;
        weight_mem[16'h257C] <= 168;
        weight_mem[16'h257D] <= 162;
        weight_mem[16'h257E] <= 161;
        weight_mem[16'h257F] <= 161;
        weight_mem[16'h2580] <= 161;
        weight_mem[16'h2581] <= 161;
        weight_mem[16'h2582] <= 161;
        weight_mem[16'h2583] <= 162;
        weight_mem[16'h2584] <= 163;
        weight_mem[16'h2585] <= 164;
        weight_mem[16'h2586] <= 170;
        weight_mem[16'h2587] <= 175;
        weight_mem[16'h2588] <= 169;
        weight_mem[16'h2589] <= 166;
        weight_mem[16'h258A] <= 170;
        weight_mem[16'h258B] <= 173;
        weight_mem[16'h258C] <= 171;
        weight_mem[16'h258D] <= 167;
        weight_mem[16'h258E] <= 171;
        weight_mem[16'h258F] <= 168;
        weight_mem[16'h2590] <= 165;
        weight_mem[16'h2591] <= 166;
        weight_mem[16'h2592] <= 168;
        weight_mem[16'h2593] <= 169;
        weight_mem[16'h2594] <= 164;
        weight_mem[16'h2595] <= 161;
        weight_mem[16'h2596] <= 161;
        weight_mem[16'h2597] <= 161;
        weight_mem[16'h2598] <= 161;
        weight_mem[16'h2599] <= 161;
        weight_mem[16'h259A] <= 161;
        weight_mem[16'h259B] <= 161;
        weight_mem[16'h259C] <= 161;
        weight_mem[16'h259D] <= 161;
        weight_mem[16'h259E] <= 162;
        weight_mem[16'h259F] <= 164;
        weight_mem[16'h25A0] <= 163;
        weight_mem[16'h25A1] <= 162;
        weight_mem[16'h25A2] <= 162;
        weight_mem[16'h25A3] <= 162;
        weight_mem[16'h25A4] <= 162;
        weight_mem[16'h25A5] <= 163;
        weight_mem[16'h25A6] <= 165;
        weight_mem[16'h25A7] <= 163;
        weight_mem[16'h25A8] <= 162;
        weight_mem[16'h25A9] <= 161;
        weight_mem[16'h25AA] <= 161;
        weight_mem[16'h25AB] <= 161;
        weight_mem[16'h25AC] <= 161;
        weight_mem[16'h25AD] <= 161;
        weight_mem[16'h25AE] <= 161;
        weight_mem[16'h25AF] <= 161;

        // layer 1 neuron 19
        weight_mem[16'h2600] <= 241;
        weight_mem[16'h2601] <= 2;
        weight_mem[16'h2602] <= 10;
        weight_mem[16'h2603] <= 253;
        weight_mem[16'h2604] <= 9;
        weight_mem[16'h2605] <= 243;
        weight_mem[16'h2606] <= 1;
        weight_mem[16'h2607] <= 244;
        weight_mem[16'h2608] <= 246;
        weight_mem[16'h2609] <= 242;
        weight_mem[16'h260A] <= 248;
        weight_mem[16'h260B] <= 242;
        weight_mem[16'h260C] <= 245;
        weight_mem[16'h260D] <= 239;
        weight_mem[16'h260E] <= 0;
        weight_mem[16'h260F] <= 252;
        weight_mem[16'h2610] <= 2;
        weight_mem[16'h2611] <= 3;
        weight_mem[16'h2612] <= 247;
        weight_mem[16'h2613] <= 6;
        weight_mem[16'h2614] <= 251;
        weight_mem[16'h2615] <= 254;
        weight_mem[16'h2616] <= 248;
        weight_mem[16'h2617] <= 246;
        weight_mem[16'h2618] <= 254;
        weight_mem[16'h2619] <= 253;
        weight_mem[16'h261A] <= 6;
        weight_mem[16'h261B] <= 2;
        weight_mem[16'h261C] <= 10;
        weight_mem[16'h261D] <= 255;
        weight_mem[16'h261E] <= 246;
        weight_mem[16'h261F] <= 254;
        weight_mem[16'h2620] <= 8;
        weight_mem[16'h2621] <= 3;
        weight_mem[16'h2622] <= 4;
        weight_mem[16'h2623] <= 247;
        weight_mem[16'h2624] <= 7;
        weight_mem[16'h2625] <= 247;
        weight_mem[16'h2626] <= 246;
        weight_mem[16'h2627] <= 242;
        weight_mem[16'h2628] <= 233;
        weight_mem[16'h2629] <= 251;
        weight_mem[16'h262A] <= 234;
        weight_mem[16'h262B] <= 253;
        weight_mem[16'h262C] <= 2;
        weight_mem[16'h262D] <= 7;
        weight_mem[16'h262E] <= 253;
        weight_mem[16'h262F] <= 247;
        weight_mem[16'h2630] <= 254;
        weight_mem[16'h2631] <= 9;
        weight_mem[16'h2632] <= 242;
        weight_mem[16'h2633] <= 245;
        weight_mem[16'h2634] <= 255;
        weight_mem[16'h2635] <= 0;
        weight_mem[16'h2636] <= 12;
        weight_mem[16'h2637] <= 18;
        weight_mem[16'h2638] <= 12;
        weight_mem[16'h2639] <= 24;
        weight_mem[16'h263A] <= 36;
        weight_mem[16'h263B] <= 43;
        weight_mem[16'h263C] <= 35;
        weight_mem[16'h263D] <= 18;
        weight_mem[16'h263E] <= 253;
        weight_mem[16'h263F] <= 245;
        weight_mem[16'h2640] <= 237;
        weight_mem[16'h2641] <= 226;
        weight_mem[16'h2642] <= 241;
        weight_mem[16'h2643] <= 243;
        weight_mem[16'h2644] <= 247;
        weight_mem[16'h2645] <= 253;
        weight_mem[16'h2646] <= 241;
        weight_mem[16'h2647] <= 239;
        weight_mem[16'h2648] <= 247;
        weight_mem[16'h2649] <= 240;
        weight_mem[16'h264A] <= 251;
        weight_mem[16'h264B] <= 3;
        weight_mem[16'h264C] <= 3;
        weight_mem[16'h264D] <= 16;
        weight_mem[16'h264E] <= 39;
        weight_mem[16'h264F] <= 20;
        weight_mem[16'h2650] <= 22;
        weight_mem[16'h2651] <= 4;
        weight_mem[16'h2652] <= 31;
        weight_mem[16'h2653] <= 28;
        weight_mem[16'h2654] <= 38;
        weight_mem[16'h2655] <= 6;
        weight_mem[16'h2656] <= 7;
        weight_mem[16'h2657] <= 238;
        weight_mem[16'h2658] <= 244;
        weight_mem[16'h2659] <= 229;
        weight_mem[16'h265A] <= 233;
        weight_mem[16'h265B] <= 208;
        weight_mem[16'h265C] <= 207;
        weight_mem[16'h265D] <= 244;
        weight_mem[16'h265E] <= 0;
        weight_mem[16'h265F] <= 250;
        weight_mem[16'h2660] <= 240;
        weight_mem[16'h2661] <= 246;
        weight_mem[16'h2662] <= 252;
        weight_mem[16'h2663] <= 17;
        weight_mem[16'h2664] <= 18;
        weight_mem[16'h2665] <= 35;
        weight_mem[16'h2666] <= 28;
        weight_mem[16'h2667] <= 7;
        weight_mem[16'h2668] <= 247;
        weight_mem[16'h2669] <= 4;
        weight_mem[16'h266A] <= 11;
        weight_mem[16'h266B] <= 41;
        weight_mem[16'h266C] <= 34;
        weight_mem[16'h266D] <= 39;
        weight_mem[16'h266E] <= 45;
        weight_mem[16'h266F] <= 37;
        weight_mem[16'h2670] <= 14;
        weight_mem[16'h2671] <= 5;
        weight_mem[16'h2672] <= 234;
        weight_mem[16'h2673] <= 206;
        weight_mem[16'h2674] <= 182;
        weight_mem[16'h2675] <= 229;
        weight_mem[16'h2676] <= 243;
        weight_mem[16'h2677] <= 0;
        weight_mem[16'h2678] <= 3;
        weight_mem[16'h2679] <= 8;
        weight_mem[16'h267A] <= 5;
        weight_mem[16'h267B] <= 31;
        weight_mem[16'h267C] <= 45;
        weight_mem[16'h267D] <= 38;
        weight_mem[16'h267E] <= 31;
        weight_mem[16'h267F] <= 5;
        weight_mem[16'h2680] <= 251;
        weight_mem[16'h2681] <= 17;
        weight_mem[16'h2682] <= 44;
        weight_mem[16'h2683] <= 90;
        weight_mem[16'h2684] <= 100;
        weight_mem[16'h2685] <= 83;
        weight_mem[16'h2686] <= 47;
        weight_mem[16'h2687] <= 35;
        weight_mem[16'h2688] <= 34;
        weight_mem[16'h2689] <= 26;
        weight_mem[16'h268A] <= 3;
        weight_mem[16'h268B] <= 228;
        weight_mem[16'h268C] <= 188;
        weight_mem[16'h268D] <= 198;
        weight_mem[16'h268E] <= 249;
        weight_mem[16'h268F] <= 242;
        weight_mem[16'h2690] <= 242;
        weight_mem[16'h2691] <= 241;
        weight_mem[16'h2692] <= 250;
        weight_mem[16'h2693] <= 32;
        weight_mem[16'h2694] <= 39;
        weight_mem[16'h2695] <= 48;
        weight_mem[16'h2696] <= 1;
        weight_mem[16'h2697] <= 1;
        weight_mem[16'h2698] <= 245;
        weight_mem[16'h2699] <= 14;
        weight_mem[16'h269A] <= 9;
        weight_mem[16'h269B] <= 30;
        weight_mem[16'h269C] <= 109;
        weight_mem[16'h269D] <= 88;
        weight_mem[16'h269E] <= 21;
        weight_mem[16'h269F] <= 17;
        weight_mem[16'h26A0] <= 9;
        weight_mem[16'h26A1] <= 38;
        weight_mem[16'h26A2] <= 19;
        weight_mem[16'h26A3] <= 245;
        weight_mem[16'h26A4] <= 213;
        weight_mem[16'h26A5] <= 219;
        weight_mem[16'h26A6] <= 236;
        weight_mem[16'h26A7] <= 10;
        weight_mem[16'h26A8] <= 2;
        weight_mem[16'h26A9] <= 252;
        weight_mem[16'h26AA] <= 0;
        weight_mem[16'h26AB] <= 29;
        weight_mem[16'h26AC] <= 48;
        weight_mem[16'h26AD] <= 15;
        weight_mem[16'h26AE] <= 253;
        weight_mem[16'h26AF] <= 247;
        weight_mem[16'h26B0] <= 247;
        weight_mem[16'h26B1] <= 220;
        weight_mem[16'h26B2] <= 189;
        weight_mem[16'h26B3] <= 203;
        weight_mem[16'h26B4] <= 38;
        weight_mem[16'h26B5] <= 29;
        weight_mem[16'h26B6] <= 0;
        weight_mem[16'h26B7] <= 9;
        weight_mem[16'h26B8] <= 43;
        weight_mem[16'h26B9] <= 69;
        weight_mem[16'h26BA] <= 58;
        weight_mem[16'h26BB] <= 3;
        weight_mem[16'h26BC] <= 255;
        weight_mem[16'h26BD] <= 4;
        weight_mem[16'h26BE] <= 252;
        weight_mem[16'h26BF] <= 248;
        weight_mem[16'h26C0] <= 2;
        weight_mem[16'h26C1] <= 7;
        weight_mem[16'h26C2] <= 1;
        weight_mem[16'h26C3] <= 5;
        weight_mem[16'h26C4] <= 21;
        weight_mem[16'h26C5] <= 234;
        weight_mem[16'h26C6] <= 221;
        weight_mem[16'h26C7] <= 242;
        weight_mem[16'h26C8] <= 242;
        weight_mem[16'h26C9] <= 177;
        weight_mem[16'h26CA] <= 128;
        weight_mem[16'h26CB] <= 181;
        weight_mem[16'h26CC] <= 16;
        weight_mem[16'h26CD] <= 1;
        weight_mem[16'h26CE] <= 242;
        weight_mem[16'h26CF] <= 253;
        weight_mem[16'h26D0] <= 12;
        weight_mem[16'h26D1] <= 43;
        weight_mem[16'h26D2] <= 10;
        weight_mem[16'h26D3] <= 243;
        weight_mem[16'h26D4] <= 247;
        weight_mem[16'h26D5] <= 12;
        weight_mem[16'h26D6] <= 5;
        weight_mem[16'h26D7] <= 1;
        weight_mem[16'h26D8] <= 10;
        weight_mem[16'h26D9] <= 248;
        weight_mem[16'h26DA] <= 7;
        weight_mem[16'h26DB] <= 254;
        weight_mem[16'h26DC] <= 6;
        weight_mem[16'h26DD] <= 250;
        weight_mem[16'h26DE] <= 242;
        weight_mem[16'h26DF] <= 238;
        weight_mem[16'h26E0] <= 218;
        weight_mem[16'h26E1] <= 167;
        weight_mem[16'h26E2] <= 161;
        weight_mem[16'h26E3] <= 244;
        weight_mem[16'h26E4] <= 8;
        weight_mem[16'h26E5] <= 228;
        weight_mem[16'h26E6] <= 242;
        weight_mem[16'h26E7] <= 245;
        weight_mem[16'h26E8] <= 0;
        weight_mem[16'h26E9] <= 246;
        weight_mem[16'h26EA] <= 10;
        weight_mem[16'h26EB] <= 230;
        weight_mem[16'h26EC] <= 233;
        weight_mem[16'h26ED] <= 255;
        weight_mem[16'h26EE] <= 9;
        weight_mem[16'h26EF] <= 12;
        weight_mem[16'h26F0] <= 254;
        weight_mem[16'h26F1] <= 11;
        weight_mem[16'h26F2] <= 9;
        weight_mem[16'h26F3] <= 12;
        weight_mem[16'h26F4] <= 22;
        weight_mem[16'h26F5] <= 249;
        weight_mem[16'h26F6] <= 2;
        weight_mem[16'h26F7] <= 240;
        weight_mem[16'h26F8] <= 244;
        weight_mem[16'h26F9] <= 222;
        weight_mem[16'h26FA] <= 2;
        weight_mem[16'h26FB] <= 38;
        weight_mem[16'h26FC] <= 251;
        weight_mem[16'h26FD] <= 255;
        weight_mem[16'h26FE] <= 7;
        weight_mem[16'h26FF] <= 4;
        weight_mem[16'h2700] <= 255;
        weight_mem[16'h2701] <= 7;
        weight_mem[16'h2702] <= 17;
        weight_mem[16'h2703] <= 12;
        weight_mem[16'h2704] <= 25;
        weight_mem[16'h2705] <= 23;
        weight_mem[16'h2706] <= 12;
        weight_mem[16'h2707] <= 4;
        weight_mem[16'h2708] <= 9;
        weight_mem[16'h2709] <= 1;
        weight_mem[16'h270A] <= 1;
        weight_mem[16'h270B] <= 16;
        weight_mem[16'h270C] <= 24;
        weight_mem[16'h270D] <= 234;
        weight_mem[16'h270E] <= 237;
        weight_mem[16'h270F] <= 241;
        weight_mem[16'h2710] <= 1;
        weight_mem[16'h2711] <= 251;
        weight_mem[16'h2712] <= 253;
        weight_mem[16'h2713] <= 14;
        weight_mem[16'h2714] <= 241;
        weight_mem[16'h2715] <= 249;
        weight_mem[16'h2716] <= 253;
        weight_mem[16'h2717] <= 246;
        weight_mem[16'h2718] <= 6;
        weight_mem[16'h2719] <= 16;
        weight_mem[16'h271A] <= 33;
        weight_mem[16'h271B] <= 33;
        weight_mem[16'h271C] <= 35;
        weight_mem[16'h271D] <= 42;
        weight_mem[16'h271E] <= 13;
        weight_mem[16'h271F] <= 252;
        weight_mem[16'h2720] <= 238;
        weight_mem[16'h2721] <= 0;
        weight_mem[16'h2722] <= 1;
        weight_mem[16'h2723] <= 32;
        weight_mem[16'h2724] <= 6;
        weight_mem[16'h2725] <= 235;
        weight_mem[16'h2726] <= 235;
        weight_mem[16'h2727] <= 213;
        weight_mem[16'h2728] <= 219;
        weight_mem[16'h2729] <= 178;
        weight_mem[16'h272A] <= 179;
        weight_mem[16'h272B] <= 193;
        weight_mem[16'h272C] <= 198;
        weight_mem[16'h272D] <= 194;
        weight_mem[16'h272E] <= 249;
        weight_mem[16'h272F] <= 237;
        weight_mem[16'h2730] <= 254;
        weight_mem[16'h2731] <= 20;
        weight_mem[16'h2732] <= 17;
        weight_mem[16'h2733] <= 12;
        weight_mem[16'h2734] <= 24;
        weight_mem[16'h2735] <= 14;
        weight_mem[16'h2736] <= 246;
        weight_mem[16'h2737] <= 8;
        weight_mem[16'h2738] <= 248;
        weight_mem[16'h2739] <= 8;
        weight_mem[16'h273A] <= 252;
        weight_mem[16'h273B] <= 18;
        weight_mem[16'h273C] <= 31;
        weight_mem[16'h273D] <= 7;
        weight_mem[16'h273E] <= 254;
        weight_mem[16'h273F] <= 247;
        weight_mem[16'h2740] <= 210;
        weight_mem[16'h2741] <= 169;
        weight_mem[16'h2742] <= 130;
        weight_mem[16'h2743] <= 147;
        weight_mem[16'h2744] <= 169;
        weight_mem[16'h2745] <= 192;
        weight_mem[16'h2746] <= 253;
        weight_mem[16'h2747] <= 4;
        weight_mem[16'h2748] <= 18;
        weight_mem[16'h2749] <= 38;
        weight_mem[16'h274A] <= 15;
        weight_mem[16'h274B] <= 14;
        weight_mem[16'h274C] <= 17;
        weight_mem[16'h274D] <= 255;
        weight_mem[16'h274E] <= 3;
        weight_mem[16'h274F] <= 244;
        weight_mem[16'h2750] <= 245;
        weight_mem[16'h2751] <= 245;
        weight_mem[16'h2752] <= 255;
        weight_mem[16'h2753] <= 12;
        weight_mem[16'h2754] <= 32;
        weight_mem[16'h2755] <= 19;
        weight_mem[16'h2756] <= 19;
        weight_mem[16'h2757] <= 10;
        weight_mem[16'h2758] <= 13;
        weight_mem[16'h2759] <= 233;
        weight_mem[16'h275A] <= 229;
        weight_mem[16'h275B] <= 209;
        weight_mem[16'h275C] <= 233;
        weight_mem[16'h275D] <= 246;
        weight_mem[16'h275E] <= 8;
        weight_mem[16'h275F] <= 9;
        weight_mem[16'h2760] <= 14;
        weight_mem[16'h2761] <= 24;
        weight_mem[16'h2762] <= 5;
        weight_mem[16'h2763] <= 3;
        weight_mem[16'h2764] <= 253;
        weight_mem[16'h2765] <= 251;
        weight_mem[16'h2766] <= 9;
        weight_mem[16'h2767] <= 242;
        weight_mem[16'h2768] <= 241;
        weight_mem[16'h2769] <= 8;
        weight_mem[16'h276A] <= 6;
        weight_mem[16'h276B] <= 251;
        weight_mem[16'h276C] <= 9;
        weight_mem[16'h276D] <= 9;
        weight_mem[16'h276E] <= 28;
        weight_mem[16'h276F] <= 1;
        weight_mem[16'h2770] <= 5;
        weight_mem[16'h2771] <= 250;
        weight_mem[16'h2772] <= 247;
        weight_mem[16'h2773] <= 241;
        weight_mem[16'h2774] <= 255;
        weight_mem[16'h2775] <= 250;
        weight_mem[16'h2776] <= 4;
        weight_mem[16'h2777] <= 11;
        weight_mem[16'h2778] <= 0;
        weight_mem[16'h2779] <= 250;
        weight_mem[16'h277A] <= 8;
        weight_mem[16'h277B] <= 3;
        weight_mem[16'h277C] <= 251;
        weight_mem[16'h277D] <= 10;
        weight_mem[16'h277E] <= 241;
        weight_mem[16'h277F] <= 9;
        weight_mem[16'h2780] <= 254;
        weight_mem[16'h2781] <= 250;
        weight_mem[16'h2782] <= 7;
        weight_mem[16'h2783] <= 250;
        weight_mem[16'h2784] <= 245;
        weight_mem[16'h2785] <= 23;
        weight_mem[16'h2786] <= 9;
        weight_mem[16'h2787] <= 24;
        weight_mem[16'h2788] <= 25;
        weight_mem[16'h2789] <= 36;
        weight_mem[16'h278A] <= 40;
        weight_mem[16'h278B] <= 33;
        weight_mem[16'h278C] <= 47;
        weight_mem[16'h278D] <= 18;
        weight_mem[16'h278E] <= 27;
        weight_mem[16'h278F] <= 13;
        weight_mem[16'h2790] <= 3;
        weight_mem[16'h2791] <= 250;
        weight_mem[16'h2792] <= 13;
        weight_mem[16'h2793] <= 5;
        weight_mem[16'h2794] <= 9;
        weight_mem[16'h2795] <= 254;
        weight_mem[16'h2796] <= 246;
        weight_mem[16'h2797] <= 10;
        weight_mem[16'h2798] <= 8;
        weight_mem[16'h2799] <= 245;
        weight_mem[16'h279A] <= 2;
        weight_mem[16'h279B] <= 1;
        weight_mem[16'h279C] <= 9;
        weight_mem[16'h279D] <= 7;
        weight_mem[16'h279E] <= 249;
        weight_mem[16'h279F] <= 11;
        weight_mem[16'h27A0] <= 251;
        weight_mem[16'h27A1] <= 252;
        weight_mem[16'h27A2] <= 255;
        weight_mem[16'h27A3] <= 15;
        weight_mem[16'h27A4] <= 2;
        weight_mem[16'h27A5] <= 22;
        weight_mem[16'h27A6] <= 255;
        weight_mem[16'h27A7] <= 4;
        weight_mem[16'h27A8] <= 253;
        weight_mem[16'h27A9] <= 9;
        weight_mem[16'h27AA] <= 252;
        weight_mem[16'h27AB] <= 238;
        weight_mem[16'h27AC] <= 10;
        weight_mem[16'h27AD] <= 244;
        weight_mem[16'h27AE] <= 254;
        weight_mem[16'h27AF] <= 250;

        // layer 1 neuron 20
        weight_mem[16'h2800] <= 0;
        weight_mem[16'h2801] <= 0;
        weight_mem[16'h2802] <= 0;
        weight_mem[16'h2803] <= 0;
        weight_mem[16'h2804] <= 0;
        weight_mem[16'h2805] <= 0;
        weight_mem[16'h2806] <= 0;
        weight_mem[16'h2807] <= 0;
        weight_mem[16'h2808] <= 0;
        weight_mem[16'h2809] <= 0;
        weight_mem[16'h280A] <= 0;
        weight_mem[16'h280B] <= 0;
        weight_mem[16'h280C] <= 0;
        weight_mem[16'h280D] <= 0;
        weight_mem[16'h280E] <= 0;
        weight_mem[16'h280F] <= 0;
        weight_mem[16'h2810] <= 0;
        weight_mem[16'h2811] <= 0;
        weight_mem[16'h2812] <= 0;
        weight_mem[16'h2813] <= 0;
        weight_mem[16'h2814] <= 0;
        weight_mem[16'h2815] <= 0;
        weight_mem[16'h2816] <= 0;
        weight_mem[16'h2817] <= 0;
        weight_mem[16'h2818] <= 0;
        weight_mem[16'h2819] <= 0;
        weight_mem[16'h281A] <= 0;
        weight_mem[16'h281B] <= 0;
        weight_mem[16'h281C] <= 0;
        weight_mem[16'h281D] <= 0;
        weight_mem[16'h281E] <= 0;
        weight_mem[16'h281F] <= 0;
        weight_mem[16'h2820] <= 0;
        weight_mem[16'h2821] <= 0;
        weight_mem[16'h2822] <= 0;
        weight_mem[16'h2823] <= 0;
        weight_mem[16'h2824] <= 0;
        weight_mem[16'h2825] <= 0;
        weight_mem[16'h2826] <= 0;
        weight_mem[16'h2827] <= 0;
        weight_mem[16'h2828] <= 0;
        weight_mem[16'h2829] <= 0;
        weight_mem[16'h282A] <= 0;
        weight_mem[16'h282B] <= 0;
        weight_mem[16'h282C] <= 0;
        weight_mem[16'h282D] <= 0;
        weight_mem[16'h282E] <= 0;
        weight_mem[16'h282F] <= 0;
        weight_mem[16'h2830] <= 0;
        weight_mem[16'h2831] <= 0;
        weight_mem[16'h2832] <= 0;
        weight_mem[16'h2833] <= 0;
        weight_mem[16'h2834] <= 0;
        weight_mem[16'h2835] <= 0;
        weight_mem[16'h2836] <= 0;
        weight_mem[16'h2837] <= 0;
        weight_mem[16'h2838] <= 0;
        weight_mem[16'h2839] <= 0;
        weight_mem[16'h283A] <= 0;
        weight_mem[16'h283B] <= 0;
        weight_mem[16'h283C] <= 0;
        weight_mem[16'h283D] <= 0;
        weight_mem[16'h283E] <= 0;
        weight_mem[16'h283F] <= 0;
        weight_mem[16'h2840] <= 0;
        weight_mem[16'h2841] <= 0;
        weight_mem[16'h2842] <= 0;
        weight_mem[16'h2843] <= 0;
        weight_mem[16'h2844] <= 0;
        weight_mem[16'h2845] <= 0;
        weight_mem[16'h2846] <= 0;
        weight_mem[16'h2847] <= 0;
        weight_mem[16'h2848] <= 0;
        weight_mem[16'h2849] <= 0;
        weight_mem[16'h284A] <= 0;
        weight_mem[16'h284B] <= 0;
        weight_mem[16'h284C] <= 0;
        weight_mem[16'h284D] <= 0;
        weight_mem[16'h284E] <= 0;
        weight_mem[16'h284F] <= 0;
        weight_mem[16'h2850] <= 0;
        weight_mem[16'h2851] <= 0;
        weight_mem[16'h2852] <= 0;
        weight_mem[16'h2853] <= 0;
        weight_mem[16'h2854] <= 0;
        weight_mem[16'h2855] <= 0;
        weight_mem[16'h2856] <= 0;
        weight_mem[16'h2857] <= 0;
        weight_mem[16'h2858] <= 0;
        weight_mem[16'h2859] <= 0;
        weight_mem[16'h285A] <= 0;
        weight_mem[16'h285B] <= 0;
        weight_mem[16'h285C] <= 0;
        weight_mem[16'h285D] <= 0;
        weight_mem[16'h285E] <= 0;
        weight_mem[16'h285F] <= 0;
        weight_mem[16'h2860] <= 0;
        weight_mem[16'h2861] <= 0;
        weight_mem[16'h2862] <= 0;
        weight_mem[16'h2863] <= 0;
        weight_mem[16'h2864] <= 0;
        weight_mem[16'h2865] <= 0;
        weight_mem[16'h2866] <= 0;
        weight_mem[16'h2867] <= 0;
        weight_mem[16'h2868] <= 0;
        weight_mem[16'h2869] <= 0;
        weight_mem[16'h286A] <= 0;
        weight_mem[16'h286B] <= 0;
        weight_mem[16'h286C] <= 0;
        weight_mem[16'h286D] <= 0;
        weight_mem[16'h286E] <= 0;
        weight_mem[16'h286F] <= 0;
        weight_mem[16'h2870] <= 0;
        weight_mem[16'h2871] <= 0;
        weight_mem[16'h2872] <= 0;
        weight_mem[16'h2873] <= 0;
        weight_mem[16'h2874] <= 0;
        weight_mem[16'h2875] <= 0;
        weight_mem[16'h2876] <= 0;
        weight_mem[16'h2877] <= 0;
        weight_mem[16'h2878] <= 0;
        weight_mem[16'h2879] <= 0;
        weight_mem[16'h287A] <= 0;
        weight_mem[16'h287B] <= 0;
        weight_mem[16'h287C] <= 0;
        weight_mem[16'h287D] <= 0;
        weight_mem[16'h287E] <= 0;
        weight_mem[16'h287F] <= 0;
        weight_mem[16'h2880] <= 0;
        weight_mem[16'h2881] <= 0;
        weight_mem[16'h2882] <= 0;
        weight_mem[16'h2883] <= 0;
        weight_mem[16'h2884] <= 0;
        weight_mem[16'h2885] <= 0;
        weight_mem[16'h2886] <= 0;
        weight_mem[16'h2887] <= 0;
        weight_mem[16'h2888] <= 0;
        weight_mem[16'h2889] <= 0;
        weight_mem[16'h288A] <= 0;
        weight_mem[16'h288B] <= 0;
        weight_mem[16'h288C] <= 0;
        weight_mem[16'h288D] <= 0;
        weight_mem[16'h288E] <= 0;
        weight_mem[16'h288F] <= 0;
        weight_mem[16'h2890] <= 0;
        weight_mem[16'h2891] <= 0;
        weight_mem[16'h2892] <= 0;
        weight_mem[16'h2893] <= 0;
        weight_mem[16'h2894] <= 0;
        weight_mem[16'h2895] <= 0;
        weight_mem[16'h2896] <= 0;
        weight_mem[16'h2897] <= 0;
        weight_mem[16'h2898] <= 0;
        weight_mem[16'h2899] <= 0;
        weight_mem[16'h289A] <= 0;
        weight_mem[16'h289B] <= 0;
        weight_mem[16'h289C] <= 0;
        weight_mem[16'h289D] <= 0;
        weight_mem[16'h289E] <= 0;
        weight_mem[16'h289F] <= 0;
        weight_mem[16'h28A0] <= 0;
        weight_mem[16'h28A1] <= 0;
        weight_mem[16'h28A2] <= 0;
        weight_mem[16'h28A3] <= 0;
        weight_mem[16'h28A4] <= 0;
        weight_mem[16'h28A5] <= 0;
        weight_mem[16'h28A6] <= 0;
        weight_mem[16'h28A7] <= 0;
        weight_mem[16'h28A8] <= 0;
        weight_mem[16'h28A9] <= 0;
        weight_mem[16'h28AA] <= 0;
        weight_mem[16'h28AB] <= 0;
        weight_mem[16'h28AC] <= 0;
        weight_mem[16'h28AD] <= 0;
        weight_mem[16'h28AE] <= 0;
        weight_mem[16'h28AF] <= 0;
        weight_mem[16'h28B0] <= 0;
        weight_mem[16'h28B1] <= 0;
        weight_mem[16'h28B2] <= 0;
        weight_mem[16'h28B3] <= 0;
        weight_mem[16'h28B4] <= 0;
        weight_mem[16'h28B5] <= 0;
        weight_mem[16'h28B6] <= 0;
        weight_mem[16'h28B7] <= 0;
        weight_mem[16'h28B8] <= 0;
        weight_mem[16'h28B9] <= 0;
        weight_mem[16'h28BA] <= 0;
        weight_mem[16'h28BB] <= 0;
        weight_mem[16'h28BC] <= 0;
        weight_mem[16'h28BD] <= 0;
        weight_mem[16'h28BE] <= 0;
        weight_mem[16'h28BF] <= 0;
        weight_mem[16'h28C0] <= 0;
        weight_mem[16'h28C1] <= 0;
        weight_mem[16'h28C2] <= 0;
        weight_mem[16'h28C3] <= 0;
        weight_mem[16'h28C4] <= 0;
        weight_mem[16'h28C5] <= 0;
        weight_mem[16'h28C6] <= 0;
        weight_mem[16'h28C7] <= 0;
        weight_mem[16'h28C8] <= 0;
        weight_mem[16'h28C9] <= 0;
        weight_mem[16'h28CA] <= 0;
        weight_mem[16'h28CB] <= 0;
        weight_mem[16'h28CC] <= 0;
        weight_mem[16'h28CD] <= 0;
        weight_mem[16'h28CE] <= 0;
        weight_mem[16'h28CF] <= 0;
        weight_mem[16'h28D0] <= 0;
        weight_mem[16'h28D1] <= 0;
        weight_mem[16'h28D2] <= 0;
        weight_mem[16'h28D3] <= 0;
        weight_mem[16'h28D4] <= 0;
        weight_mem[16'h28D5] <= 0;
        weight_mem[16'h28D6] <= 0;
        weight_mem[16'h28D7] <= 0;
        weight_mem[16'h28D8] <= 0;
        weight_mem[16'h28D9] <= 0;
        weight_mem[16'h28DA] <= 0;
        weight_mem[16'h28DB] <= 0;
        weight_mem[16'h28DC] <= 0;
        weight_mem[16'h28DD] <= 0;
        weight_mem[16'h28DE] <= 0;
        weight_mem[16'h28DF] <= 0;
        weight_mem[16'h28E0] <= 0;
        weight_mem[16'h28E1] <= 0;
        weight_mem[16'h28E2] <= 0;
        weight_mem[16'h28E3] <= 0;
        weight_mem[16'h28E4] <= 0;
        weight_mem[16'h28E5] <= 0;
        weight_mem[16'h28E6] <= 0;
        weight_mem[16'h28E7] <= 0;
        weight_mem[16'h28E8] <= 0;
        weight_mem[16'h28E9] <= 0;
        weight_mem[16'h28EA] <= 0;
        weight_mem[16'h28EB] <= 0;
        weight_mem[16'h28EC] <= 0;
        weight_mem[16'h28ED] <= 0;
        weight_mem[16'h28EE] <= 0;
        weight_mem[16'h28EF] <= 0;
        weight_mem[16'h28F0] <= 0;
        weight_mem[16'h28F1] <= 0;
        weight_mem[16'h28F2] <= 0;
        weight_mem[16'h28F3] <= 0;
        weight_mem[16'h28F4] <= 0;
        weight_mem[16'h28F5] <= 0;
        weight_mem[16'h28F6] <= 0;
        weight_mem[16'h28F7] <= 0;
        weight_mem[16'h28F8] <= 0;
        weight_mem[16'h28F9] <= 0;
        weight_mem[16'h28FA] <= 0;
        weight_mem[16'h28FB] <= 0;
        weight_mem[16'h28FC] <= 0;
        weight_mem[16'h28FD] <= 0;
        weight_mem[16'h28FE] <= 0;
        weight_mem[16'h28FF] <= 0;
        weight_mem[16'h2900] <= 0;
        weight_mem[16'h2901] <= 0;
        weight_mem[16'h2902] <= 0;
        weight_mem[16'h2903] <= 0;
        weight_mem[16'h2904] <= 0;
        weight_mem[16'h2905] <= 0;
        weight_mem[16'h2906] <= 0;
        weight_mem[16'h2907] <= 0;
        weight_mem[16'h2908] <= 0;
        weight_mem[16'h2909] <= 0;
        weight_mem[16'h290A] <= 0;
        weight_mem[16'h290B] <= 0;
        weight_mem[16'h290C] <= 0;
        weight_mem[16'h290D] <= 0;
        weight_mem[16'h290E] <= 0;
        weight_mem[16'h290F] <= 0;
        weight_mem[16'h2910] <= 0;
        weight_mem[16'h2911] <= 0;
        weight_mem[16'h2912] <= 0;
        weight_mem[16'h2913] <= 0;
        weight_mem[16'h2914] <= 0;
        weight_mem[16'h2915] <= 0;
        weight_mem[16'h2916] <= 0;
        weight_mem[16'h2917] <= 0;
        weight_mem[16'h2918] <= 0;
        weight_mem[16'h2919] <= 0;
        weight_mem[16'h291A] <= 0;
        weight_mem[16'h291B] <= 0;
        weight_mem[16'h291C] <= 0;
        weight_mem[16'h291D] <= 0;
        weight_mem[16'h291E] <= 0;
        weight_mem[16'h291F] <= 0;
        weight_mem[16'h2920] <= 0;
        weight_mem[16'h2921] <= 0;
        weight_mem[16'h2922] <= 0;
        weight_mem[16'h2923] <= 0;
        weight_mem[16'h2924] <= 0;
        weight_mem[16'h2925] <= 0;
        weight_mem[16'h2926] <= 0;
        weight_mem[16'h2927] <= 0;
        weight_mem[16'h2928] <= 0;
        weight_mem[16'h2929] <= 0;
        weight_mem[16'h292A] <= 0;
        weight_mem[16'h292B] <= 0;
        weight_mem[16'h292C] <= 0;
        weight_mem[16'h292D] <= 0;
        weight_mem[16'h292E] <= 0;
        weight_mem[16'h292F] <= 0;
        weight_mem[16'h2930] <= 0;
        weight_mem[16'h2931] <= 0;
        weight_mem[16'h2932] <= 0;
        weight_mem[16'h2933] <= 0;
        weight_mem[16'h2934] <= 0;
        weight_mem[16'h2935] <= 0;
        weight_mem[16'h2936] <= 0;
        weight_mem[16'h2937] <= 0;
        weight_mem[16'h2938] <= 0;
        weight_mem[16'h2939] <= 0;
        weight_mem[16'h293A] <= 0;
        weight_mem[16'h293B] <= 0;
        weight_mem[16'h293C] <= 0;
        weight_mem[16'h293D] <= 0;
        weight_mem[16'h293E] <= 0;
        weight_mem[16'h293F] <= 0;
        weight_mem[16'h2940] <= 0;
        weight_mem[16'h2941] <= 0;
        weight_mem[16'h2942] <= 0;
        weight_mem[16'h2943] <= 0;
        weight_mem[16'h2944] <= 0;
        weight_mem[16'h2945] <= 0;
        weight_mem[16'h2946] <= 0;
        weight_mem[16'h2947] <= 0;
        weight_mem[16'h2948] <= 0;
        weight_mem[16'h2949] <= 0;
        weight_mem[16'h294A] <= 0;
        weight_mem[16'h294B] <= 0;
        weight_mem[16'h294C] <= 0;
        weight_mem[16'h294D] <= 0;
        weight_mem[16'h294E] <= 0;
        weight_mem[16'h294F] <= 0;
        weight_mem[16'h2950] <= 0;
        weight_mem[16'h2951] <= 0;
        weight_mem[16'h2952] <= 0;
        weight_mem[16'h2953] <= 0;
        weight_mem[16'h2954] <= 0;
        weight_mem[16'h2955] <= 0;
        weight_mem[16'h2956] <= 0;
        weight_mem[16'h2957] <= 0;
        weight_mem[16'h2958] <= 0;
        weight_mem[16'h2959] <= 0;
        weight_mem[16'h295A] <= 0;
        weight_mem[16'h295B] <= 0;
        weight_mem[16'h295C] <= 0;
        weight_mem[16'h295D] <= 0;
        weight_mem[16'h295E] <= 0;
        weight_mem[16'h295F] <= 0;
        weight_mem[16'h2960] <= 0;
        weight_mem[16'h2961] <= 0;
        weight_mem[16'h2962] <= 0;
        weight_mem[16'h2963] <= 0;
        weight_mem[16'h2964] <= 0;
        weight_mem[16'h2965] <= 0;
        weight_mem[16'h2966] <= 0;
        weight_mem[16'h2967] <= 0;
        weight_mem[16'h2968] <= 0;
        weight_mem[16'h2969] <= 0;
        weight_mem[16'h296A] <= 0;
        weight_mem[16'h296B] <= 0;
        weight_mem[16'h296C] <= 0;
        weight_mem[16'h296D] <= 0;
        weight_mem[16'h296E] <= 0;
        weight_mem[16'h296F] <= 0;
        weight_mem[16'h2970] <= 0;
        weight_mem[16'h2971] <= 0;
        weight_mem[16'h2972] <= 0;
        weight_mem[16'h2973] <= 0;
        weight_mem[16'h2974] <= 0;
        weight_mem[16'h2975] <= 0;
        weight_mem[16'h2976] <= 0;
        weight_mem[16'h2977] <= 0;
        weight_mem[16'h2978] <= 0;
        weight_mem[16'h2979] <= 0;
        weight_mem[16'h297A] <= 0;
        weight_mem[16'h297B] <= 0;
        weight_mem[16'h297C] <= 0;
        weight_mem[16'h297D] <= 0;
        weight_mem[16'h297E] <= 0;
        weight_mem[16'h297F] <= 0;
        weight_mem[16'h2980] <= 0;
        weight_mem[16'h2981] <= 0;
        weight_mem[16'h2982] <= 0;
        weight_mem[16'h2983] <= 0;
        weight_mem[16'h2984] <= 0;
        weight_mem[16'h2985] <= 0;
        weight_mem[16'h2986] <= 0;
        weight_mem[16'h2987] <= 0;
        weight_mem[16'h2988] <= 0;
        weight_mem[16'h2989] <= 0;
        weight_mem[16'h298A] <= 0;
        weight_mem[16'h298B] <= 0;
        weight_mem[16'h298C] <= 0;
        weight_mem[16'h298D] <= 0;
        weight_mem[16'h298E] <= 0;
        weight_mem[16'h298F] <= 0;
        weight_mem[16'h2990] <= 0;
        weight_mem[16'h2991] <= 0;
        weight_mem[16'h2992] <= 0;
        weight_mem[16'h2993] <= 0;
        weight_mem[16'h2994] <= 0;
        weight_mem[16'h2995] <= 0;
        weight_mem[16'h2996] <= 0;
        weight_mem[16'h2997] <= 0;
        weight_mem[16'h2998] <= 0;
        weight_mem[16'h2999] <= 0;
        weight_mem[16'h299A] <= 0;
        weight_mem[16'h299B] <= 0;
        weight_mem[16'h299C] <= 0;
        weight_mem[16'h299D] <= 0;
        weight_mem[16'h299E] <= 0;
        weight_mem[16'h299F] <= 0;
        weight_mem[16'h29A0] <= 0;
        weight_mem[16'h29A1] <= 0;
        weight_mem[16'h29A2] <= 0;
        weight_mem[16'h29A3] <= 0;
        weight_mem[16'h29A4] <= 0;
        weight_mem[16'h29A5] <= 0;
        weight_mem[16'h29A6] <= 0;
        weight_mem[16'h29A7] <= 0;
        weight_mem[16'h29A8] <= 0;
        weight_mem[16'h29A9] <= 0;
        weight_mem[16'h29AA] <= 0;
        weight_mem[16'h29AB] <= 0;
        weight_mem[16'h29AC] <= 0;
        weight_mem[16'h29AD] <= 0;
        weight_mem[16'h29AE] <= 0;
        weight_mem[16'h29AF] <= 0;

        // layer 1 neuron 21
        weight_mem[16'h2A00] <= 177;
        weight_mem[16'h2A01] <= 177;
        weight_mem[16'h2A02] <= 177;
        weight_mem[16'h2A03] <= 177;
        weight_mem[16'h2A04] <= 177;
        weight_mem[16'h2A05] <= 177;
        weight_mem[16'h2A06] <= 177;
        weight_mem[16'h2A07] <= 177;
        weight_mem[16'h2A08] <= 177;
        weight_mem[16'h2A09] <= 177;
        weight_mem[16'h2A0A] <= 177;
        weight_mem[16'h2A0B] <= 177;
        weight_mem[16'h2A0C] <= 177;
        weight_mem[16'h2A0D] <= 177;
        weight_mem[16'h2A0E] <= 177;
        weight_mem[16'h2A0F] <= 177;
        weight_mem[16'h2A10] <= 177;
        weight_mem[16'h2A11] <= 178;
        weight_mem[16'h2A12] <= 183;
        weight_mem[16'h2A13] <= 179;
        weight_mem[16'h2A14] <= 177;
        weight_mem[16'h2A15] <= 177;
        weight_mem[16'h2A16] <= 177;
        weight_mem[16'h2A17] <= 177;
        weight_mem[16'h2A18] <= 177;
        weight_mem[16'h2A19] <= 177;
        weight_mem[16'h2A1A] <= 177;
        weight_mem[16'h2A1B] <= 177;
        weight_mem[16'h2A1C] <= 177;
        weight_mem[16'h2A1D] <= 177;
        weight_mem[16'h2A1E] <= 177;
        weight_mem[16'h2A1F] <= 177;
        weight_mem[16'h2A20] <= 176;
        weight_mem[16'h2A21] <= 177;
        weight_mem[16'h2A22] <= 178;
        weight_mem[16'h2A23] <= 177;
        weight_mem[16'h2A24] <= 177;
        weight_mem[16'h2A25] <= 179;
        weight_mem[16'h2A26] <= 179;
        weight_mem[16'h2A27] <= 178;
        weight_mem[16'h2A28] <= 179;
        weight_mem[16'h2A29] <= 187;
        weight_mem[16'h2A2A] <= 193;
        weight_mem[16'h2A2B] <= 186;
        weight_mem[16'h2A2C] <= 177;
        weight_mem[16'h2A2D] <= 177;
        weight_mem[16'h2A2E] <= 177;
        weight_mem[16'h2A2F] <= 177;
        weight_mem[16'h2A30] <= 177;
        weight_mem[16'h2A31] <= 177;
        weight_mem[16'h2A32] <= 177;
        weight_mem[16'h2A33] <= 177;
        weight_mem[16'h2A34] <= 177;
        weight_mem[16'h2A35] <= 177;
        weight_mem[16'h2A36] <= 178;
        weight_mem[16'h2A37] <= 177;
        weight_mem[16'h2A38] <= 170;
        weight_mem[16'h2A39] <= 165;
        weight_mem[16'h2A3A] <= 167;
        weight_mem[16'h2A3B] <= 170;
        weight_mem[16'h2A3C] <= 173;
        weight_mem[16'h2A3D] <= 181;
        weight_mem[16'h2A3E] <= 182;
        weight_mem[16'h2A3F] <= 187;
        weight_mem[16'h2A40] <= 202;
        weight_mem[16'h2A41] <= 208;
        weight_mem[16'h2A42] <= 202;
        weight_mem[16'h2A43] <= 190;
        weight_mem[16'h2A44] <= 179;
        weight_mem[16'h2A45] <= 177;
        weight_mem[16'h2A46] <= 177;
        weight_mem[16'h2A47] <= 177;
        weight_mem[16'h2A48] <= 177;
        weight_mem[16'h2A49] <= 177;
        weight_mem[16'h2A4A] <= 176;
        weight_mem[16'h2A4B] <= 175;
        weight_mem[16'h2A4C] <= 177;
        weight_mem[16'h2A4D] <= 183;
        weight_mem[16'h2A4E] <= 197;
        weight_mem[16'h2A4F] <= 220;
        weight_mem[16'h2A50] <= 224;
        weight_mem[16'h2A51] <= 215;
        weight_mem[16'h2A52] <= 196;
        weight_mem[16'h2A53] <= 181;
        weight_mem[16'h2A54] <= 186;
        weight_mem[16'h2A55] <= 195;
        weight_mem[16'h2A56] <= 215;
        weight_mem[16'h2A57] <= 232;
        weight_mem[16'h2A58] <= 242;
        weight_mem[16'h2A59] <= 239;
        weight_mem[16'h2A5A] <= 226;
        weight_mem[16'h2A5B] <= 202;
        weight_mem[16'h2A5C] <= 181;
        weight_mem[16'h2A5D] <= 177;
        weight_mem[16'h2A5E] <= 177;
        weight_mem[16'h2A5F] <= 177;
        weight_mem[16'h2A60] <= 177;
        weight_mem[16'h2A61] <= 176;
        weight_mem[16'h2A62] <= 167;
        weight_mem[16'h2A63] <= 159;
        weight_mem[16'h2A64] <= 172;
        weight_mem[16'h2A65] <= 179;
        weight_mem[16'h2A66] <= 170;
        weight_mem[16'h2A67] <= 211;
        weight_mem[16'h2A68] <= 217;
        weight_mem[16'h2A69] <= 219;
        weight_mem[16'h2A6A] <= 217;
        weight_mem[16'h2A6B] <= 222;
        weight_mem[16'h2A6C] <= 230;
        weight_mem[16'h2A6D] <= 239;
        weight_mem[16'h2A6E] <= 245;
        weight_mem[16'h2A6F] <= 246;
        weight_mem[16'h2A70] <= 249;
        weight_mem[16'h2A71] <= 250;
        weight_mem[16'h2A72] <= 234;
        weight_mem[16'h2A73] <= 199;
        weight_mem[16'h2A74] <= 180;
        weight_mem[16'h2A75] <= 182;
        weight_mem[16'h2A76] <= 178;
        weight_mem[16'h2A77] <= 177;
        weight_mem[16'h2A78] <= 173;
        weight_mem[16'h2A79] <= 155;
        weight_mem[16'h2A7A] <= 158;
        weight_mem[16'h2A7B] <= 162;
        weight_mem[16'h2A7C] <= 175;
        weight_mem[16'h2A7D] <= 173;
        weight_mem[16'h2A7E] <= 131;
        weight_mem[16'h2A7F] <= 176;
        weight_mem[16'h2A80] <= 196;
        weight_mem[16'h2A81] <= 222;
        weight_mem[16'h2A82] <= 249;
        weight_mem[16'h2A83] <= 0;
        weight_mem[16'h2A84] <= 0;
        weight_mem[16'h2A85] <= 0;
        weight_mem[16'h2A86] <= 0;
        weight_mem[16'h2A87] <= 252;
        weight_mem[16'h2A88] <= 250;
        weight_mem[16'h2A89] <= 248;
        weight_mem[16'h2A8A] <= 222;
        weight_mem[16'h2A8B] <= 196;
        weight_mem[16'h2A8C] <= 183;
        weight_mem[16'h2A8D] <= 181;
        weight_mem[16'h2A8E] <= 178;
        weight_mem[16'h2A8F] <= 178;
        weight_mem[16'h2A90] <= 171;
        weight_mem[16'h2A91] <= 139;
        weight_mem[16'h2A92] <= 139;
        weight_mem[16'h2A93] <= 146;
        weight_mem[16'h2A94] <= 171;
        weight_mem[16'h2A95] <= 187;
        weight_mem[16'h2A96] <= 181;
        weight_mem[16'h2A97] <= 253;
        weight_mem[16'h2A98] <= 0;
        weight_mem[16'h2A99] <= 0;
        weight_mem[16'h2A9A] <= 255;
        weight_mem[16'h2A9B] <= 250;
        weight_mem[16'h2A9C] <= 255;
        weight_mem[16'h2A9D] <= 0;
        weight_mem[16'h2A9E] <= 0;
        weight_mem[16'h2A9F] <= 0;
        weight_mem[16'h2AA0] <= 235;
        weight_mem[16'h2AA1] <= 219;
        weight_mem[16'h2AA2] <= 205;
        weight_mem[16'h2AA3] <= 189;
        weight_mem[16'h2AA4] <= 173;
        weight_mem[16'h2AA5] <= 177;
        weight_mem[16'h2AA6] <= 177;
        weight_mem[16'h2AA7] <= 177;
        weight_mem[16'h2AA8] <= 174;
        weight_mem[16'h2AA9] <= 155;
        weight_mem[16'h2AAA] <= 141;
        weight_mem[16'h2AAB] <= 144;
        weight_mem[16'h2AAC] <= 150;
        weight_mem[16'h2AAD] <= 167;
        weight_mem[16'h2AAE] <= 225;
        weight_mem[16'h2AAF] <= 254;
        weight_mem[16'h2AB0] <= 250;
        weight_mem[16'h2AB1] <= 244;
        weight_mem[16'h2AB2] <= 254;
        weight_mem[16'h2AB3] <= 255;
        weight_mem[16'h2AB4] <= 255;
        weight_mem[16'h2AB5] <= 252;
        weight_mem[16'h2AB6] <= 0;
        weight_mem[16'h2AB7] <= 0;
        weight_mem[16'h2AB8] <= 234;
        weight_mem[16'h2AB9] <= 207;
        weight_mem[16'h2ABA] <= 212;
        weight_mem[16'h2ABB] <= 191;
        weight_mem[16'h2ABC] <= 175;
        weight_mem[16'h2ABD] <= 177;
        weight_mem[16'h2ABE] <= 177;
        weight_mem[16'h2ABF] <= 177;
        weight_mem[16'h2AC0] <= 177;
        weight_mem[16'h2AC1] <= 173;
        weight_mem[16'h2AC2] <= 169;
        weight_mem[16'h2AC3] <= 168;
        weight_mem[16'h2AC4] <= 160;
        weight_mem[16'h2AC5] <= 181;
        weight_mem[16'h2AC6] <= 242;
        weight_mem[16'h2AC7] <= 249;
        weight_mem[16'h2AC8] <= 249;
        weight_mem[16'h2AC9] <= 245;
        weight_mem[16'h2ACA] <= 249;
        weight_mem[16'h2ACB] <= 244;
        weight_mem[16'h2ACC] <= 227;
        weight_mem[16'h2ACD] <= 250;
        weight_mem[16'h2ACE] <= 0;
        weight_mem[16'h2ACF] <= 255;
        weight_mem[16'h2AD0] <= 233;
        weight_mem[16'h2AD1] <= 220;
        weight_mem[16'h2AD2] <= 219;
        weight_mem[16'h2AD3] <= 187;
        weight_mem[16'h2AD4] <= 176;
        weight_mem[16'h2AD5] <= 178;
        weight_mem[16'h2AD6] <= 177;
        weight_mem[16'h2AD7] <= 177;
        weight_mem[16'h2AD8] <= 177;
        weight_mem[16'h2AD9] <= 177;
        weight_mem[16'h2ADA] <= 180;
        weight_mem[16'h2ADB] <= 186;
        weight_mem[16'h2ADC] <= 195;
        weight_mem[16'h2ADD] <= 199;
        weight_mem[16'h2ADE] <= 217;
        weight_mem[16'h2ADF] <= 221;
        weight_mem[16'h2AE0] <= 243;
        weight_mem[16'h2AE1] <= 251;
        weight_mem[16'h2AE2] <= 248;
        weight_mem[16'h2AE3] <= 239;
        weight_mem[16'h2AE4] <= 225;
        weight_mem[16'h2AE5] <= 249;
        weight_mem[16'h2AE6] <= 0;
        weight_mem[16'h2AE7] <= 239;
        weight_mem[16'h2AE8] <= 207;
        weight_mem[16'h2AE9] <= 228;
        weight_mem[16'h2AEA] <= 224;
        weight_mem[16'h2AEB] <= 186;
        weight_mem[16'h2AEC] <= 182;
        weight_mem[16'h2AED] <= 177;
        weight_mem[16'h2AEE] <= 175;
        weight_mem[16'h2AEF] <= 175;
        weight_mem[16'h2AF0] <= 177;
        weight_mem[16'h2AF1] <= 177;
        weight_mem[16'h2AF2] <= 179;
        weight_mem[16'h2AF3] <= 193;
        weight_mem[16'h2AF4] <= 213;
        weight_mem[16'h2AF5] <= 212;
        weight_mem[16'h2AF6] <= 202;
        weight_mem[16'h2AF7] <= 209;
        weight_mem[16'h2AF8] <= 249;
        weight_mem[16'h2AF9] <= 254;
        weight_mem[16'h2AFA] <= 251;
        weight_mem[16'h2AFB] <= 244;
        weight_mem[16'h2AFC] <= 244;
        weight_mem[16'h2AFD] <= 254;
        weight_mem[16'h2AFE] <= 255;
        weight_mem[16'h2AFF] <= 209;
        weight_mem[16'h2B00] <= 184;
        weight_mem[16'h2B01] <= 206;
        weight_mem[16'h2B02] <= 203;
        weight_mem[16'h2B03] <= 172;
        weight_mem[16'h2B04] <= 169;
        weight_mem[16'h2B05] <= 164;
        weight_mem[16'h2B06] <= 162;
        weight_mem[16'h2B07] <= 167;
        weight_mem[16'h2B08] <= 177;
        weight_mem[16'h2B09] <= 177;
        weight_mem[16'h2B0A] <= 183;
        weight_mem[16'h2B0B] <= 197;
        weight_mem[16'h2B0C] <= 209;
        weight_mem[16'h2B0D] <= 208;
        weight_mem[16'h2B0E] <= 213;
        weight_mem[16'h2B0F] <= 208;
        weight_mem[16'h2B10] <= 234;
        weight_mem[16'h2B11] <= 245;
        weight_mem[16'h2B12] <= 241;
        weight_mem[16'h2B13] <= 234;
        weight_mem[16'h2B14] <= 248;
        weight_mem[16'h2B15] <= 255;
        weight_mem[16'h2B16] <= 254;
        weight_mem[16'h2B17] <= 214;
        weight_mem[16'h2B18] <= 205;
        weight_mem[16'h2B19] <= 202;
        weight_mem[16'h2B1A] <= 181;
        weight_mem[16'h2B1B] <= 152;
        weight_mem[16'h2B1C] <= 169;
        weight_mem[16'h2B1D] <= 170;
        weight_mem[16'h2B1E] <= 174;
        weight_mem[16'h2B1F] <= 176;
        weight_mem[16'h2B20] <= 177;
        weight_mem[16'h2B21] <= 177;
        weight_mem[16'h2B22] <= 184;
        weight_mem[16'h2B23] <= 195;
        weight_mem[16'h2B24] <= 203;
        weight_mem[16'h2B25] <= 214;
        weight_mem[16'h2B26] <= 229;
        weight_mem[16'h2B27] <= 227;
        weight_mem[16'h2B28] <= 225;
        weight_mem[16'h2B29] <= 225;
        weight_mem[16'h2B2A] <= 221;
        weight_mem[16'h2B2B] <= 232;
        weight_mem[16'h2B2C] <= 250;
        weight_mem[16'h2B2D] <= 0;
        weight_mem[16'h2B2E] <= 252;
        weight_mem[16'h2B2F] <= 202;
        weight_mem[16'h2B30] <= 208;
        weight_mem[16'h2B31] <= 217;
        weight_mem[16'h2B32] <= 209;
        weight_mem[16'h2B33] <= 178;
        weight_mem[16'h2B34] <= 176;
        weight_mem[16'h2B35] <= 176;
        weight_mem[16'h2B36] <= 177;
        weight_mem[16'h2B37] <= 177;
        weight_mem[16'h2B38] <= 177;
        weight_mem[16'h2B39] <= 177;
        weight_mem[16'h2B3A] <= 178;
        weight_mem[16'h2B3B] <= 184;
        weight_mem[16'h2B3C] <= 193;
        weight_mem[16'h2B3D] <= 218;
        weight_mem[16'h2B3E] <= 236;
        weight_mem[16'h2B3F] <= 243;
        weight_mem[16'h2B40] <= 245;
        weight_mem[16'h2B41] <= 244;
        weight_mem[16'h2B42] <= 241;
        weight_mem[16'h2B43] <= 241;
        weight_mem[16'h2B44] <= 236;
        weight_mem[16'h2B45] <= 247;
        weight_mem[16'h2B46] <= 239;
        weight_mem[16'h2B47] <= 175;
        weight_mem[16'h2B48] <= 176;
        weight_mem[16'h2B49] <= 196;
        weight_mem[16'h2B4A] <= 202;
        weight_mem[16'h2B4B] <= 196;
        weight_mem[16'h2B4C] <= 179;
        weight_mem[16'h2B4D] <= 175;
        weight_mem[16'h2B4E] <= 177;
        weight_mem[16'h2B4F] <= 177;
        weight_mem[16'h2B50] <= 177;
        weight_mem[16'h2B51] <= 177;
        weight_mem[16'h2B52] <= 176;
        weight_mem[16'h2B53] <= 176;
        weight_mem[16'h2B54] <= 184;
        weight_mem[16'h2B55] <= 207;
        weight_mem[16'h2B56] <= 213;
        weight_mem[16'h2B57] <= 221;
        weight_mem[16'h2B58] <= 237;
        weight_mem[16'h2B59] <= 242;
        weight_mem[16'h2B5A] <= 243;
        weight_mem[16'h2B5B] <= 247;
        weight_mem[16'h2B5C] <= 233;
        weight_mem[16'h2B5D] <= 251;
        weight_mem[16'h2B5E] <= 252;
        weight_mem[16'h2B5F] <= 220;
        weight_mem[16'h2B60] <= 212;
        weight_mem[16'h2B61] <= 205;
        weight_mem[16'h2B62] <= 200;
        weight_mem[16'h2B63] <= 185;
        weight_mem[16'h2B64] <= 177;
        weight_mem[16'h2B65] <= 177;
        weight_mem[16'h2B66] <= 177;
        weight_mem[16'h2B67] <= 177;
        weight_mem[16'h2B68] <= 177;
        weight_mem[16'h2B69] <= 177;
        weight_mem[16'h2B6A] <= 177;
        weight_mem[16'h2B6B] <= 177;
        weight_mem[16'h2B6C] <= 178;
        weight_mem[16'h2B6D] <= 186;
        weight_mem[16'h2B6E] <= 180;
        weight_mem[16'h2B6F] <= 186;
        weight_mem[16'h2B70] <= 217;
        weight_mem[16'h2B71] <= 224;
        weight_mem[16'h2B72] <= 231;
        weight_mem[16'h2B73] <= 240;
        weight_mem[16'h2B74] <= 226;
        weight_mem[16'h2B75] <= 251;
        weight_mem[16'h2B76] <= 248;
        weight_mem[16'h2B77] <= 163;
        weight_mem[16'h2B78] <= 158;
        weight_mem[16'h2B79] <= 185;
        weight_mem[16'h2B7A] <= 184;
        weight_mem[16'h2B7B] <= 175;
        weight_mem[16'h2B7C] <= 176;
        weight_mem[16'h2B7D] <= 177;
        weight_mem[16'h2B7E] <= 177;
        weight_mem[16'h2B7F] <= 177;
        weight_mem[16'h2B80] <= 177;
        weight_mem[16'h2B81] <= 177;
        weight_mem[16'h2B82] <= 177;
        weight_mem[16'h2B83] <= 177;
        weight_mem[16'h2B84] <= 177;
        weight_mem[16'h2B85] <= 176;
        weight_mem[16'h2B86] <= 173;
        weight_mem[16'h2B87] <= 175;
        weight_mem[16'h2B88] <= 186;
        weight_mem[16'h2B89] <= 188;
        weight_mem[16'h2B8A] <= 194;
        weight_mem[16'h2B8B] <= 203;
        weight_mem[16'h2B8C] <= 194;
        weight_mem[16'h2B8D] <= 239;
        weight_mem[16'h2B8E] <= 214;
        weight_mem[16'h2B8F] <= 128;
        weight_mem[16'h2B90] <= 139;
        weight_mem[16'h2B91] <= 178;
        weight_mem[16'h2B92] <= 184;
        weight_mem[16'h2B93] <= 178;
        weight_mem[16'h2B94] <= 177;
        weight_mem[16'h2B95] <= 177;
        weight_mem[16'h2B96] <= 177;
        weight_mem[16'h2B97] <= 177;
        weight_mem[16'h2B98] <= 177;
        weight_mem[16'h2B99] <= 177;
        weight_mem[16'h2B9A] <= 177;
        weight_mem[16'h2B9B] <= 177;
        weight_mem[16'h2B9C] <= 177;
        weight_mem[16'h2B9D] <= 177;
        weight_mem[16'h2B9E] <= 176;
        weight_mem[16'h2B9F] <= 178;
        weight_mem[16'h2BA0] <= 180;
        weight_mem[16'h2BA1] <= 178;
        weight_mem[16'h2BA2] <= 177;
        weight_mem[16'h2BA3] <= 184;
        weight_mem[16'h2BA4] <= 198;
        weight_mem[16'h2BA5] <= 239;
        weight_mem[16'h2BA6] <= 202;
        weight_mem[16'h2BA7] <= 171;
        weight_mem[16'h2BA8] <= 168;
        weight_mem[16'h2BA9] <= 176;
        weight_mem[16'h2BAA] <= 178;
        weight_mem[16'h2BAB] <= 177;
        weight_mem[16'h2BAC] <= 177;
        weight_mem[16'h2BAD] <= 177;
        weight_mem[16'h2BAE] <= 177;
        weight_mem[16'h2BAF] <= 177;

        // layer 1 neuron 22
        weight_mem[16'h2C00] <= 0;
        weight_mem[16'h2C01] <= 0;
        weight_mem[16'h2C02] <= 0;
        weight_mem[16'h2C03] <= 0;
        weight_mem[16'h2C04] <= 0;
        weight_mem[16'h2C05] <= 0;
        weight_mem[16'h2C06] <= 0;
        weight_mem[16'h2C07] <= 0;
        weight_mem[16'h2C08] <= 0;
        weight_mem[16'h2C09] <= 0;
        weight_mem[16'h2C0A] <= 0;
        weight_mem[16'h2C0B] <= 0;
        weight_mem[16'h2C0C] <= 0;
        weight_mem[16'h2C0D] <= 0;
        weight_mem[16'h2C0E] <= 0;
        weight_mem[16'h2C0F] <= 0;
        weight_mem[16'h2C10] <= 0;
        weight_mem[16'h2C11] <= 0;
        weight_mem[16'h2C12] <= 0;
        weight_mem[16'h2C13] <= 0;
        weight_mem[16'h2C14] <= 0;
        weight_mem[16'h2C15] <= 0;
        weight_mem[16'h2C16] <= 0;
        weight_mem[16'h2C17] <= 0;
        weight_mem[16'h2C18] <= 0;
        weight_mem[16'h2C19] <= 0;
        weight_mem[16'h2C1A] <= 0;
        weight_mem[16'h2C1B] <= 0;
        weight_mem[16'h2C1C] <= 0;
        weight_mem[16'h2C1D] <= 0;
        weight_mem[16'h2C1E] <= 0;
        weight_mem[16'h2C1F] <= 0;
        weight_mem[16'h2C20] <= 0;
        weight_mem[16'h2C21] <= 0;
        weight_mem[16'h2C22] <= 0;
        weight_mem[16'h2C23] <= 0;
        weight_mem[16'h2C24] <= 0;
        weight_mem[16'h2C25] <= 0;
        weight_mem[16'h2C26] <= 0;
        weight_mem[16'h2C27] <= 0;
        weight_mem[16'h2C28] <= 0;
        weight_mem[16'h2C29] <= 0;
        weight_mem[16'h2C2A] <= 0;
        weight_mem[16'h2C2B] <= 0;
        weight_mem[16'h2C2C] <= 0;
        weight_mem[16'h2C2D] <= 0;
        weight_mem[16'h2C2E] <= 0;
        weight_mem[16'h2C2F] <= 0;
        weight_mem[16'h2C30] <= 0;
        weight_mem[16'h2C31] <= 0;
        weight_mem[16'h2C32] <= 0;
        weight_mem[16'h2C33] <= 0;
        weight_mem[16'h2C34] <= 0;
        weight_mem[16'h2C35] <= 0;
        weight_mem[16'h2C36] <= 0;
        weight_mem[16'h2C37] <= 0;
        weight_mem[16'h2C38] <= 0;
        weight_mem[16'h2C39] <= 0;
        weight_mem[16'h2C3A] <= 0;
        weight_mem[16'h2C3B] <= 0;
        weight_mem[16'h2C3C] <= 0;
        weight_mem[16'h2C3D] <= 0;
        weight_mem[16'h2C3E] <= 0;
        weight_mem[16'h2C3F] <= 0;
        weight_mem[16'h2C40] <= 0;
        weight_mem[16'h2C41] <= 0;
        weight_mem[16'h2C42] <= 0;
        weight_mem[16'h2C43] <= 0;
        weight_mem[16'h2C44] <= 0;
        weight_mem[16'h2C45] <= 0;
        weight_mem[16'h2C46] <= 0;
        weight_mem[16'h2C47] <= 0;
        weight_mem[16'h2C48] <= 0;
        weight_mem[16'h2C49] <= 0;
        weight_mem[16'h2C4A] <= 0;
        weight_mem[16'h2C4B] <= 0;
        weight_mem[16'h2C4C] <= 0;
        weight_mem[16'h2C4D] <= 0;
        weight_mem[16'h2C4E] <= 0;
        weight_mem[16'h2C4F] <= 0;
        weight_mem[16'h2C50] <= 0;
        weight_mem[16'h2C51] <= 0;
        weight_mem[16'h2C52] <= 0;
        weight_mem[16'h2C53] <= 0;
        weight_mem[16'h2C54] <= 0;
        weight_mem[16'h2C55] <= 0;
        weight_mem[16'h2C56] <= 0;
        weight_mem[16'h2C57] <= 0;
        weight_mem[16'h2C58] <= 0;
        weight_mem[16'h2C59] <= 0;
        weight_mem[16'h2C5A] <= 0;
        weight_mem[16'h2C5B] <= 0;
        weight_mem[16'h2C5C] <= 0;
        weight_mem[16'h2C5D] <= 0;
        weight_mem[16'h2C5E] <= 0;
        weight_mem[16'h2C5F] <= 0;
        weight_mem[16'h2C60] <= 0;
        weight_mem[16'h2C61] <= 0;
        weight_mem[16'h2C62] <= 0;
        weight_mem[16'h2C63] <= 0;
        weight_mem[16'h2C64] <= 0;
        weight_mem[16'h2C65] <= 0;
        weight_mem[16'h2C66] <= 0;
        weight_mem[16'h2C67] <= 0;
        weight_mem[16'h2C68] <= 0;
        weight_mem[16'h2C69] <= 0;
        weight_mem[16'h2C6A] <= 0;
        weight_mem[16'h2C6B] <= 0;
        weight_mem[16'h2C6C] <= 0;
        weight_mem[16'h2C6D] <= 0;
        weight_mem[16'h2C6E] <= 0;
        weight_mem[16'h2C6F] <= 0;
        weight_mem[16'h2C70] <= 0;
        weight_mem[16'h2C71] <= 0;
        weight_mem[16'h2C72] <= 0;
        weight_mem[16'h2C73] <= 0;
        weight_mem[16'h2C74] <= 0;
        weight_mem[16'h2C75] <= 0;
        weight_mem[16'h2C76] <= 0;
        weight_mem[16'h2C77] <= 0;
        weight_mem[16'h2C78] <= 0;
        weight_mem[16'h2C79] <= 0;
        weight_mem[16'h2C7A] <= 0;
        weight_mem[16'h2C7B] <= 0;
        weight_mem[16'h2C7C] <= 0;
        weight_mem[16'h2C7D] <= 0;
        weight_mem[16'h2C7E] <= 0;
        weight_mem[16'h2C7F] <= 0;
        weight_mem[16'h2C80] <= 0;
        weight_mem[16'h2C81] <= 0;
        weight_mem[16'h2C82] <= 0;
        weight_mem[16'h2C83] <= 0;
        weight_mem[16'h2C84] <= 0;
        weight_mem[16'h2C85] <= 0;
        weight_mem[16'h2C86] <= 0;
        weight_mem[16'h2C87] <= 0;
        weight_mem[16'h2C88] <= 0;
        weight_mem[16'h2C89] <= 0;
        weight_mem[16'h2C8A] <= 0;
        weight_mem[16'h2C8B] <= 0;
        weight_mem[16'h2C8C] <= 0;
        weight_mem[16'h2C8D] <= 0;
        weight_mem[16'h2C8E] <= 0;
        weight_mem[16'h2C8F] <= 0;
        weight_mem[16'h2C90] <= 0;
        weight_mem[16'h2C91] <= 0;
        weight_mem[16'h2C92] <= 0;
        weight_mem[16'h2C93] <= 0;
        weight_mem[16'h2C94] <= 0;
        weight_mem[16'h2C95] <= 0;
        weight_mem[16'h2C96] <= 0;
        weight_mem[16'h2C97] <= 0;
        weight_mem[16'h2C98] <= 0;
        weight_mem[16'h2C99] <= 0;
        weight_mem[16'h2C9A] <= 0;
        weight_mem[16'h2C9B] <= 0;
        weight_mem[16'h2C9C] <= 0;
        weight_mem[16'h2C9D] <= 0;
        weight_mem[16'h2C9E] <= 0;
        weight_mem[16'h2C9F] <= 0;
        weight_mem[16'h2CA0] <= 0;
        weight_mem[16'h2CA1] <= 0;
        weight_mem[16'h2CA2] <= 0;
        weight_mem[16'h2CA3] <= 0;
        weight_mem[16'h2CA4] <= 0;
        weight_mem[16'h2CA5] <= 0;
        weight_mem[16'h2CA6] <= 0;
        weight_mem[16'h2CA7] <= 0;
        weight_mem[16'h2CA8] <= 0;
        weight_mem[16'h2CA9] <= 0;
        weight_mem[16'h2CAA] <= 0;
        weight_mem[16'h2CAB] <= 0;
        weight_mem[16'h2CAC] <= 0;
        weight_mem[16'h2CAD] <= 0;
        weight_mem[16'h2CAE] <= 0;
        weight_mem[16'h2CAF] <= 0;
        weight_mem[16'h2CB0] <= 0;
        weight_mem[16'h2CB1] <= 0;
        weight_mem[16'h2CB2] <= 0;
        weight_mem[16'h2CB3] <= 0;
        weight_mem[16'h2CB4] <= 0;
        weight_mem[16'h2CB5] <= 0;
        weight_mem[16'h2CB6] <= 0;
        weight_mem[16'h2CB7] <= 0;
        weight_mem[16'h2CB8] <= 0;
        weight_mem[16'h2CB9] <= 0;
        weight_mem[16'h2CBA] <= 0;
        weight_mem[16'h2CBB] <= 0;
        weight_mem[16'h2CBC] <= 0;
        weight_mem[16'h2CBD] <= 0;
        weight_mem[16'h2CBE] <= 0;
        weight_mem[16'h2CBF] <= 0;
        weight_mem[16'h2CC0] <= 0;
        weight_mem[16'h2CC1] <= 0;
        weight_mem[16'h2CC2] <= 0;
        weight_mem[16'h2CC3] <= 0;
        weight_mem[16'h2CC4] <= 0;
        weight_mem[16'h2CC5] <= 0;
        weight_mem[16'h2CC6] <= 0;
        weight_mem[16'h2CC7] <= 0;
        weight_mem[16'h2CC8] <= 0;
        weight_mem[16'h2CC9] <= 0;
        weight_mem[16'h2CCA] <= 0;
        weight_mem[16'h2CCB] <= 0;
        weight_mem[16'h2CCC] <= 0;
        weight_mem[16'h2CCD] <= 0;
        weight_mem[16'h2CCE] <= 0;
        weight_mem[16'h2CCF] <= 0;
        weight_mem[16'h2CD0] <= 0;
        weight_mem[16'h2CD1] <= 0;
        weight_mem[16'h2CD2] <= 0;
        weight_mem[16'h2CD3] <= 0;
        weight_mem[16'h2CD4] <= 0;
        weight_mem[16'h2CD5] <= 0;
        weight_mem[16'h2CD6] <= 0;
        weight_mem[16'h2CD7] <= 0;
        weight_mem[16'h2CD8] <= 0;
        weight_mem[16'h2CD9] <= 0;
        weight_mem[16'h2CDA] <= 0;
        weight_mem[16'h2CDB] <= 0;
        weight_mem[16'h2CDC] <= 0;
        weight_mem[16'h2CDD] <= 0;
        weight_mem[16'h2CDE] <= 0;
        weight_mem[16'h2CDF] <= 0;
        weight_mem[16'h2CE0] <= 0;
        weight_mem[16'h2CE1] <= 0;
        weight_mem[16'h2CE2] <= 0;
        weight_mem[16'h2CE3] <= 0;
        weight_mem[16'h2CE4] <= 0;
        weight_mem[16'h2CE5] <= 0;
        weight_mem[16'h2CE6] <= 0;
        weight_mem[16'h2CE7] <= 0;
        weight_mem[16'h2CE8] <= 0;
        weight_mem[16'h2CE9] <= 0;
        weight_mem[16'h2CEA] <= 0;
        weight_mem[16'h2CEB] <= 0;
        weight_mem[16'h2CEC] <= 0;
        weight_mem[16'h2CED] <= 0;
        weight_mem[16'h2CEE] <= 0;
        weight_mem[16'h2CEF] <= 0;
        weight_mem[16'h2CF0] <= 0;
        weight_mem[16'h2CF1] <= 0;
        weight_mem[16'h2CF2] <= 0;
        weight_mem[16'h2CF3] <= 0;
        weight_mem[16'h2CF4] <= 0;
        weight_mem[16'h2CF5] <= 0;
        weight_mem[16'h2CF6] <= 0;
        weight_mem[16'h2CF7] <= 0;
        weight_mem[16'h2CF8] <= 0;
        weight_mem[16'h2CF9] <= 0;
        weight_mem[16'h2CFA] <= 0;
        weight_mem[16'h2CFB] <= 0;
        weight_mem[16'h2CFC] <= 0;
        weight_mem[16'h2CFD] <= 0;
        weight_mem[16'h2CFE] <= 0;
        weight_mem[16'h2CFF] <= 0;
        weight_mem[16'h2D00] <= 0;
        weight_mem[16'h2D01] <= 0;
        weight_mem[16'h2D02] <= 0;
        weight_mem[16'h2D03] <= 0;
        weight_mem[16'h2D04] <= 0;
        weight_mem[16'h2D05] <= 0;
        weight_mem[16'h2D06] <= 0;
        weight_mem[16'h2D07] <= 0;
        weight_mem[16'h2D08] <= 0;
        weight_mem[16'h2D09] <= 0;
        weight_mem[16'h2D0A] <= 0;
        weight_mem[16'h2D0B] <= 0;
        weight_mem[16'h2D0C] <= 0;
        weight_mem[16'h2D0D] <= 0;
        weight_mem[16'h2D0E] <= 0;
        weight_mem[16'h2D0F] <= 0;
        weight_mem[16'h2D10] <= 0;
        weight_mem[16'h2D11] <= 0;
        weight_mem[16'h2D12] <= 0;
        weight_mem[16'h2D13] <= 0;
        weight_mem[16'h2D14] <= 0;
        weight_mem[16'h2D15] <= 0;
        weight_mem[16'h2D16] <= 0;
        weight_mem[16'h2D17] <= 0;
        weight_mem[16'h2D18] <= 0;
        weight_mem[16'h2D19] <= 0;
        weight_mem[16'h2D1A] <= 0;
        weight_mem[16'h2D1B] <= 0;
        weight_mem[16'h2D1C] <= 0;
        weight_mem[16'h2D1D] <= 0;
        weight_mem[16'h2D1E] <= 0;
        weight_mem[16'h2D1F] <= 0;
        weight_mem[16'h2D20] <= 0;
        weight_mem[16'h2D21] <= 0;
        weight_mem[16'h2D22] <= 0;
        weight_mem[16'h2D23] <= 0;
        weight_mem[16'h2D24] <= 0;
        weight_mem[16'h2D25] <= 0;
        weight_mem[16'h2D26] <= 0;
        weight_mem[16'h2D27] <= 0;
        weight_mem[16'h2D28] <= 0;
        weight_mem[16'h2D29] <= 0;
        weight_mem[16'h2D2A] <= 0;
        weight_mem[16'h2D2B] <= 0;
        weight_mem[16'h2D2C] <= 0;
        weight_mem[16'h2D2D] <= 0;
        weight_mem[16'h2D2E] <= 0;
        weight_mem[16'h2D2F] <= 0;
        weight_mem[16'h2D30] <= 0;
        weight_mem[16'h2D31] <= 0;
        weight_mem[16'h2D32] <= 0;
        weight_mem[16'h2D33] <= 0;
        weight_mem[16'h2D34] <= 0;
        weight_mem[16'h2D35] <= 0;
        weight_mem[16'h2D36] <= 0;
        weight_mem[16'h2D37] <= 0;
        weight_mem[16'h2D38] <= 0;
        weight_mem[16'h2D39] <= 0;
        weight_mem[16'h2D3A] <= 0;
        weight_mem[16'h2D3B] <= 0;
        weight_mem[16'h2D3C] <= 0;
        weight_mem[16'h2D3D] <= 0;
        weight_mem[16'h2D3E] <= 0;
        weight_mem[16'h2D3F] <= 0;
        weight_mem[16'h2D40] <= 0;
        weight_mem[16'h2D41] <= 0;
        weight_mem[16'h2D42] <= 0;
        weight_mem[16'h2D43] <= 0;
        weight_mem[16'h2D44] <= 0;
        weight_mem[16'h2D45] <= 0;
        weight_mem[16'h2D46] <= 0;
        weight_mem[16'h2D47] <= 0;
        weight_mem[16'h2D48] <= 0;
        weight_mem[16'h2D49] <= 0;
        weight_mem[16'h2D4A] <= 0;
        weight_mem[16'h2D4B] <= 0;
        weight_mem[16'h2D4C] <= 0;
        weight_mem[16'h2D4D] <= 0;
        weight_mem[16'h2D4E] <= 0;
        weight_mem[16'h2D4F] <= 0;
        weight_mem[16'h2D50] <= 0;
        weight_mem[16'h2D51] <= 0;
        weight_mem[16'h2D52] <= 0;
        weight_mem[16'h2D53] <= 0;
        weight_mem[16'h2D54] <= 0;
        weight_mem[16'h2D55] <= 0;
        weight_mem[16'h2D56] <= 0;
        weight_mem[16'h2D57] <= 0;
        weight_mem[16'h2D58] <= 0;
        weight_mem[16'h2D59] <= 0;
        weight_mem[16'h2D5A] <= 0;
        weight_mem[16'h2D5B] <= 0;
        weight_mem[16'h2D5C] <= 0;
        weight_mem[16'h2D5D] <= 0;
        weight_mem[16'h2D5E] <= 0;
        weight_mem[16'h2D5F] <= 0;
        weight_mem[16'h2D60] <= 0;
        weight_mem[16'h2D61] <= 0;
        weight_mem[16'h2D62] <= 0;
        weight_mem[16'h2D63] <= 0;
        weight_mem[16'h2D64] <= 0;
        weight_mem[16'h2D65] <= 0;
        weight_mem[16'h2D66] <= 0;
        weight_mem[16'h2D67] <= 0;
        weight_mem[16'h2D68] <= 0;
        weight_mem[16'h2D69] <= 0;
        weight_mem[16'h2D6A] <= 0;
        weight_mem[16'h2D6B] <= 0;
        weight_mem[16'h2D6C] <= 0;
        weight_mem[16'h2D6D] <= 0;
        weight_mem[16'h2D6E] <= 0;
        weight_mem[16'h2D6F] <= 0;
        weight_mem[16'h2D70] <= 0;
        weight_mem[16'h2D71] <= 0;
        weight_mem[16'h2D72] <= 0;
        weight_mem[16'h2D73] <= 0;
        weight_mem[16'h2D74] <= 0;
        weight_mem[16'h2D75] <= 0;
        weight_mem[16'h2D76] <= 0;
        weight_mem[16'h2D77] <= 0;
        weight_mem[16'h2D78] <= 0;
        weight_mem[16'h2D79] <= 0;
        weight_mem[16'h2D7A] <= 0;
        weight_mem[16'h2D7B] <= 0;
        weight_mem[16'h2D7C] <= 0;
        weight_mem[16'h2D7D] <= 0;
        weight_mem[16'h2D7E] <= 0;
        weight_mem[16'h2D7F] <= 0;
        weight_mem[16'h2D80] <= 0;
        weight_mem[16'h2D81] <= 0;
        weight_mem[16'h2D82] <= 0;
        weight_mem[16'h2D83] <= 0;
        weight_mem[16'h2D84] <= 0;
        weight_mem[16'h2D85] <= 0;
        weight_mem[16'h2D86] <= 0;
        weight_mem[16'h2D87] <= 0;
        weight_mem[16'h2D88] <= 0;
        weight_mem[16'h2D89] <= 0;
        weight_mem[16'h2D8A] <= 0;
        weight_mem[16'h2D8B] <= 0;
        weight_mem[16'h2D8C] <= 0;
        weight_mem[16'h2D8D] <= 0;
        weight_mem[16'h2D8E] <= 0;
        weight_mem[16'h2D8F] <= 0;
        weight_mem[16'h2D90] <= 0;
        weight_mem[16'h2D91] <= 0;
        weight_mem[16'h2D92] <= 0;
        weight_mem[16'h2D93] <= 0;
        weight_mem[16'h2D94] <= 0;
        weight_mem[16'h2D95] <= 0;
        weight_mem[16'h2D96] <= 0;
        weight_mem[16'h2D97] <= 0;
        weight_mem[16'h2D98] <= 0;
        weight_mem[16'h2D99] <= 0;
        weight_mem[16'h2D9A] <= 0;
        weight_mem[16'h2D9B] <= 0;
        weight_mem[16'h2D9C] <= 0;
        weight_mem[16'h2D9D] <= 0;
        weight_mem[16'h2D9E] <= 0;
        weight_mem[16'h2D9F] <= 0;
        weight_mem[16'h2DA0] <= 0;
        weight_mem[16'h2DA1] <= 0;
        weight_mem[16'h2DA2] <= 0;
        weight_mem[16'h2DA3] <= 0;
        weight_mem[16'h2DA4] <= 0;
        weight_mem[16'h2DA5] <= 0;
        weight_mem[16'h2DA6] <= 0;
        weight_mem[16'h2DA7] <= 0;
        weight_mem[16'h2DA8] <= 0;
        weight_mem[16'h2DA9] <= 0;
        weight_mem[16'h2DAA] <= 0;
        weight_mem[16'h2DAB] <= 0;
        weight_mem[16'h2DAC] <= 0;
        weight_mem[16'h2DAD] <= 0;
        weight_mem[16'h2DAE] <= 0;
        weight_mem[16'h2DAF] <= 0;

        // layer 1 neuron 23
        weight_mem[16'h2E00] <= 0;
        weight_mem[16'h2E01] <= 0;
        weight_mem[16'h2E02] <= 0;
        weight_mem[16'h2E03] <= 0;
        weight_mem[16'h2E04] <= 0;
        weight_mem[16'h2E05] <= 0;
        weight_mem[16'h2E06] <= 0;
        weight_mem[16'h2E07] <= 0;
        weight_mem[16'h2E08] <= 0;
        weight_mem[16'h2E09] <= 0;
        weight_mem[16'h2E0A] <= 0;
        weight_mem[16'h2E0B] <= 0;
        weight_mem[16'h2E0C] <= 0;
        weight_mem[16'h2E0D] <= 0;
        weight_mem[16'h2E0E] <= 0;
        weight_mem[16'h2E0F] <= 0;
        weight_mem[16'h2E10] <= 0;
        weight_mem[16'h2E11] <= 0;
        weight_mem[16'h2E12] <= 0;
        weight_mem[16'h2E13] <= 0;
        weight_mem[16'h2E14] <= 0;
        weight_mem[16'h2E15] <= 0;
        weight_mem[16'h2E16] <= 0;
        weight_mem[16'h2E17] <= 0;
        weight_mem[16'h2E18] <= 0;
        weight_mem[16'h2E19] <= 0;
        weight_mem[16'h2E1A] <= 0;
        weight_mem[16'h2E1B] <= 0;
        weight_mem[16'h2E1C] <= 0;
        weight_mem[16'h2E1D] <= 0;
        weight_mem[16'h2E1E] <= 0;
        weight_mem[16'h2E1F] <= 0;
        weight_mem[16'h2E20] <= 0;
        weight_mem[16'h2E21] <= 0;
        weight_mem[16'h2E22] <= 0;
        weight_mem[16'h2E23] <= 0;
        weight_mem[16'h2E24] <= 0;
        weight_mem[16'h2E25] <= 0;
        weight_mem[16'h2E26] <= 0;
        weight_mem[16'h2E27] <= 0;
        weight_mem[16'h2E28] <= 0;
        weight_mem[16'h2E29] <= 0;
        weight_mem[16'h2E2A] <= 0;
        weight_mem[16'h2E2B] <= 0;
        weight_mem[16'h2E2C] <= 0;
        weight_mem[16'h2E2D] <= 0;
        weight_mem[16'h2E2E] <= 0;
        weight_mem[16'h2E2F] <= 0;
        weight_mem[16'h2E30] <= 0;
        weight_mem[16'h2E31] <= 0;
        weight_mem[16'h2E32] <= 0;
        weight_mem[16'h2E33] <= 0;
        weight_mem[16'h2E34] <= 0;
        weight_mem[16'h2E35] <= 0;
        weight_mem[16'h2E36] <= 0;
        weight_mem[16'h2E37] <= 0;
        weight_mem[16'h2E38] <= 0;
        weight_mem[16'h2E39] <= 0;
        weight_mem[16'h2E3A] <= 0;
        weight_mem[16'h2E3B] <= 0;
        weight_mem[16'h2E3C] <= 0;
        weight_mem[16'h2E3D] <= 0;
        weight_mem[16'h2E3E] <= 0;
        weight_mem[16'h2E3F] <= 0;
        weight_mem[16'h2E40] <= 0;
        weight_mem[16'h2E41] <= 0;
        weight_mem[16'h2E42] <= 0;
        weight_mem[16'h2E43] <= 0;
        weight_mem[16'h2E44] <= 0;
        weight_mem[16'h2E45] <= 0;
        weight_mem[16'h2E46] <= 0;
        weight_mem[16'h2E47] <= 0;
        weight_mem[16'h2E48] <= 0;
        weight_mem[16'h2E49] <= 0;
        weight_mem[16'h2E4A] <= 0;
        weight_mem[16'h2E4B] <= 0;
        weight_mem[16'h2E4C] <= 0;
        weight_mem[16'h2E4D] <= 0;
        weight_mem[16'h2E4E] <= 0;
        weight_mem[16'h2E4F] <= 0;
        weight_mem[16'h2E50] <= 0;
        weight_mem[16'h2E51] <= 0;
        weight_mem[16'h2E52] <= 0;
        weight_mem[16'h2E53] <= 0;
        weight_mem[16'h2E54] <= 0;
        weight_mem[16'h2E55] <= 0;
        weight_mem[16'h2E56] <= 0;
        weight_mem[16'h2E57] <= 0;
        weight_mem[16'h2E58] <= 0;
        weight_mem[16'h2E59] <= 0;
        weight_mem[16'h2E5A] <= 0;
        weight_mem[16'h2E5B] <= 0;
        weight_mem[16'h2E5C] <= 0;
        weight_mem[16'h2E5D] <= 0;
        weight_mem[16'h2E5E] <= 0;
        weight_mem[16'h2E5F] <= 0;
        weight_mem[16'h2E60] <= 0;
        weight_mem[16'h2E61] <= 0;
        weight_mem[16'h2E62] <= 0;
        weight_mem[16'h2E63] <= 0;
        weight_mem[16'h2E64] <= 0;
        weight_mem[16'h2E65] <= 0;
        weight_mem[16'h2E66] <= 0;
        weight_mem[16'h2E67] <= 0;
        weight_mem[16'h2E68] <= 0;
        weight_mem[16'h2E69] <= 0;
        weight_mem[16'h2E6A] <= 0;
        weight_mem[16'h2E6B] <= 0;
        weight_mem[16'h2E6C] <= 0;
        weight_mem[16'h2E6D] <= 0;
        weight_mem[16'h2E6E] <= 0;
        weight_mem[16'h2E6F] <= 0;
        weight_mem[16'h2E70] <= 0;
        weight_mem[16'h2E71] <= 0;
        weight_mem[16'h2E72] <= 0;
        weight_mem[16'h2E73] <= 0;
        weight_mem[16'h2E74] <= 0;
        weight_mem[16'h2E75] <= 0;
        weight_mem[16'h2E76] <= 0;
        weight_mem[16'h2E77] <= 0;
        weight_mem[16'h2E78] <= 0;
        weight_mem[16'h2E79] <= 0;
        weight_mem[16'h2E7A] <= 0;
        weight_mem[16'h2E7B] <= 0;
        weight_mem[16'h2E7C] <= 0;
        weight_mem[16'h2E7D] <= 0;
        weight_mem[16'h2E7E] <= 0;
        weight_mem[16'h2E7F] <= 0;
        weight_mem[16'h2E80] <= 0;
        weight_mem[16'h2E81] <= 0;
        weight_mem[16'h2E82] <= 0;
        weight_mem[16'h2E83] <= 0;
        weight_mem[16'h2E84] <= 0;
        weight_mem[16'h2E85] <= 0;
        weight_mem[16'h2E86] <= 0;
        weight_mem[16'h2E87] <= 0;
        weight_mem[16'h2E88] <= 0;
        weight_mem[16'h2E89] <= 0;
        weight_mem[16'h2E8A] <= 0;
        weight_mem[16'h2E8B] <= 0;
        weight_mem[16'h2E8C] <= 0;
        weight_mem[16'h2E8D] <= 0;
        weight_mem[16'h2E8E] <= 0;
        weight_mem[16'h2E8F] <= 0;
        weight_mem[16'h2E90] <= 0;
        weight_mem[16'h2E91] <= 0;
        weight_mem[16'h2E92] <= 0;
        weight_mem[16'h2E93] <= 0;
        weight_mem[16'h2E94] <= 0;
        weight_mem[16'h2E95] <= 0;
        weight_mem[16'h2E96] <= 0;
        weight_mem[16'h2E97] <= 0;
        weight_mem[16'h2E98] <= 0;
        weight_mem[16'h2E99] <= 0;
        weight_mem[16'h2E9A] <= 0;
        weight_mem[16'h2E9B] <= 0;
        weight_mem[16'h2E9C] <= 0;
        weight_mem[16'h2E9D] <= 0;
        weight_mem[16'h2E9E] <= 0;
        weight_mem[16'h2E9F] <= 0;
        weight_mem[16'h2EA0] <= 0;
        weight_mem[16'h2EA1] <= 0;
        weight_mem[16'h2EA2] <= 0;
        weight_mem[16'h2EA3] <= 0;
        weight_mem[16'h2EA4] <= 0;
        weight_mem[16'h2EA5] <= 0;
        weight_mem[16'h2EA6] <= 0;
        weight_mem[16'h2EA7] <= 0;
        weight_mem[16'h2EA8] <= 0;
        weight_mem[16'h2EA9] <= 0;
        weight_mem[16'h2EAA] <= 0;
        weight_mem[16'h2EAB] <= 0;
        weight_mem[16'h2EAC] <= 0;
        weight_mem[16'h2EAD] <= 0;
        weight_mem[16'h2EAE] <= 0;
        weight_mem[16'h2EAF] <= 0;
        weight_mem[16'h2EB0] <= 0;
        weight_mem[16'h2EB1] <= 0;
        weight_mem[16'h2EB2] <= 0;
        weight_mem[16'h2EB3] <= 0;
        weight_mem[16'h2EB4] <= 0;
        weight_mem[16'h2EB5] <= 0;
        weight_mem[16'h2EB6] <= 0;
        weight_mem[16'h2EB7] <= 0;
        weight_mem[16'h2EB8] <= 0;
        weight_mem[16'h2EB9] <= 0;
        weight_mem[16'h2EBA] <= 0;
        weight_mem[16'h2EBB] <= 0;
        weight_mem[16'h2EBC] <= 0;
        weight_mem[16'h2EBD] <= 0;
        weight_mem[16'h2EBE] <= 0;
        weight_mem[16'h2EBF] <= 0;
        weight_mem[16'h2EC0] <= 0;
        weight_mem[16'h2EC1] <= 0;
        weight_mem[16'h2EC2] <= 0;
        weight_mem[16'h2EC3] <= 0;
        weight_mem[16'h2EC4] <= 0;
        weight_mem[16'h2EC5] <= 0;
        weight_mem[16'h2EC6] <= 0;
        weight_mem[16'h2EC7] <= 0;
        weight_mem[16'h2EC8] <= 0;
        weight_mem[16'h2EC9] <= 0;
        weight_mem[16'h2ECA] <= 0;
        weight_mem[16'h2ECB] <= 0;
        weight_mem[16'h2ECC] <= 0;
        weight_mem[16'h2ECD] <= 0;
        weight_mem[16'h2ECE] <= 0;
        weight_mem[16'h2ECF] <= 0;
        weight_mem[16'h2ED0] <= 0;
        weight_mem[16'h2ED1] <= 0;
        weight_mem[16'h2ED2] <= 0;
        weight_mem[16'h2ED3] <= 0;
        weight_mem[16'h2ED4] <= 0;
        weight_mem[16'h2ED5] <= 0;
        weight_mem[16'h2ED6] <= 0;
        weight_mem[16'h2ED7] <= 0;
        weight_mem[16'h2ED8] <= 0;
        weight_mem[16'h2ED9] <= 0;
        weight_mem[16'h2EDA] <= 0;
        weight_mem[16'h2EDB] <= 0;
        weight_mem[16'h2EDC] <= 0;
        weight_mem[16'h2EDD] <= 0;
        weight_mem[16'h2EDE] <= 0;
        weight_mem[16'h2EDF] <= 0;
        weight_mem[16'h2EE0] <= 0;
        weight_mem[16'h2EE1] <= 0;
        weight_mem[16'h2EE2] <= 0;
        weight_mem[16'h2EE3] <= 0;
        weight_mem[16'h2EE4] <= 0;
        weight_mem[16'h2EE5] <= 0;
        weight_mem[16'h2EE6] <= 0;
        weight_mem[16'h2EE7] <= 0;
        weight_mem[16'h2EE8] <= 0;
        weight_mem[16'h2EE9] <= 0;
        weight_mem[16'h2EEA] <= 0;
        weight_mem[16'h2EEB] <= 0;
        weight_mem[16'h2EEC] <= 0;
        weight_mem[16'h2EED] <= 0;
        weight_mem[16'h2EEE] <= 0;
        weight_mem[16'h2EEF] <= 0;
        weight_mem[16'h2EF0] <= 0;
        weight_mem[16'h2EF1] <= 0;
        weight_mem[16'h2EF2] <= 0;
        weight_mem[16'h2EF3] <= 0;
        weight_mem[16'h2EF4] <= 0;
        weight_mem[16'h2EF5] <= 0;
        weight_mem[16'h2EF6] <= 0;
        weight_mem[16'h2EF7] <= 0;
        weight_mem[16'h2EF8] <= 0;
        weight_mem[16'h2EF9] <= 0;
        weight_mem[16'h2EFA] <= 0;
        weight_mem[16'h2EFB] <= 0;
        weight_mem[16'h2EFC] <= 0;
        weight_mem[16'h2EFD] <= 0;
        weight_mem[16'h2EFE] <= 0;
        weight_mem[16'h2EFF] <= 0;
        weight_mem[16'h2F00] <= 0;
        weight_mem[16'h2F01] <= 0;
        weight_mem[16'h2F02] <= 0;
        weight_mem[16'h2F03] <= 0;
        weight_mem[16'h2F04] <= 0;
        weight_mem[16'h2F05] <= 0;
        weight_mem[16'h2F06] <= 0;
        weight_mem[16'h2F07] <= 0;
        weight_mem[16'h2F08] <= 0;
        weight_mem[16'h2F09] <= 0;
        weight_mem[16'h2F0A] <= 0;
        weight_mem[16'h2F0B] <= 0;
        weight_mem[16'h2F0C] <= 0;
        weight_mem[16'h2F0D] <= 0;
        weight_mem[16'h2F0E] <= 0;
        weight_mem[16'h2F0F] <= 0;
        weight_mem[16'h2F10] <= 0;
        weight_mem[16'h2F11] <= 0;
        weight_mem[16'h2F12] <= 0;
        weight_mem[16'h2F13] <= 0;
        weight_mem[16'h2F14] <= 0;
        weight_mem[16'h2F15] <= 0;
        weight_mem[16'h2F16] <= 0;
        weight_mem[16'h2F17] <= 0;
        weight_mem[16'h2F18] <= 0;
        weight_mem[16'h2F19] <= 0;
        weight_mem[16'h2F1A] <= 0;
        weight_mem[16'h2F1B] <= 0;
        weight_mem[16'h2F1C] <= 0;
        weight_mem[16'h2F1D] <= 0;
        weight_mem[16'h2F1E] <= 0;
        weight_mem[16'h2F1F] <= 0;
        weight_mem[16'h2F20] <= 0;
        weight_mem[16'h2F21] <= 0;
        weight_mem[16'h2F22] <= 0;
        weight_mem[16'h2F23] <= 0;
        weight_mem[16'h2F24] <= 0;
        weight_mem[16'h2F25] <= 0;
        weight_mem[16'h2F26] <= 0;
        weight_mem[16'h2F27] <= 0;
        weight_mem[16'h2F28] <= 0;
        weight_mem[16'h2F29] <= 0;
        weight_mem[16'h2F2A] <= 0;
        weight_mem[16'h2F2B] <= 0;
        weight_mem[16'h2F2C] <= 0;
        weight_mem[16'h2F2D] <= 0;
        weight_mem[16'h2F2E] <= 0;
        weight_mem[16'h2F2F] <= 0;
        weight_mem[16'h2F30] <= 0;
        weight_mem[16'h2F31] <= 0;
        weight_mem[16'h2F32] <= 0;
        weight_mem[16'h2F33] <= 0;
        weight_mem[16'h2F34] <= 0;
        weight_mem[16'h2F35] <= 0;
        weight_mem[16'h2F36] <= 0;
        weight_mem[16'h2F37] <= 0;
        weight_mem[16'h2F38] <= 0;
        weight_mem[16'h2F39] <= 0;
        weight_mem[16'h2F3A] <= 0;
        weight_mem[16'h2F3B] <= 0;
        weight_mem[16'h2F3C] <= 0;
        weight_mem[16'h2F3D] <= 0;
        weight_mem[16'h2F3E] <= 0;
        weight_mem[16'h2F3F] <= 0;
        weight_mem[16'h2F40] <= 0;
        weight_mem[16'h2F41] <= 0;
        weight_mem[16'h2F42] <= 0;
        weight_mem[16'h2F43] <= 0;
        weight_mem[16'h2F44] <= 0;
        weight_mem[16'h2F45] <= 0;
        weight_mem[16'h2F46] <= 0;
        weight_mem[16'h2F47] <= 0;
        weight_mem[16'h2F48] <= 0;
        weight_mem[16'h2F49] <= 0;
        weight_mem[16'h2F4A] <= 0;
        weight_mem[16'h2F4B] <= 0;
        weight_mem[16'h2F4C] <= 0;
        weight_mem[16'h2F4D] <= 0;
        weight_mem[16'h2F4E] <= 0;
        weight_mem[16'h2F4F] <= 0;
        weight_mem[16'h2F50] <= 0;
        weight_mem[16'h2F51] <= 0;
        weight_mem[16'h2F52] <= 0;
        weight_mem[16'h2F53] <= 0;
        weight_mem[16'h2F54] <= 0;
        weight_mem[16'h2F55] <= 0;
        weight_mem[16'h2F56] <= 0;
        weight_mem[16'h2F57] <= 0;
        weight_mem[16'h2F58] <= 0;
        weight_mem[16'h2F59] <= 0;
        weight_mem[16'h2F5A] <= 0;
        weight_mem[16'h2F5B] <= 0;
        weight_mem[16'h2F5C] <= 0;
        weight_mem[16'h2F5D] <= 0;
        weight_mem[16'h2F5E] <= 0;
        weight_mem[16'h2F5F] <= 0;
        weight_mem[16'h2F60] <= 0;
        weight_mem[16'h2F61] <= 0;
        weight_mem[16'h2F62] <= 0;
        weight_mem[16'h2F63] <= 0;
        weight_mem[16'h2F64] <= 0;
        weight_mem[16'h2F65] <= 0;
        weight_mem[16'h2F66] <= 0;
        weight_mem[16'h2F67] <= 0;
        weight_mem[16'h2F68] <= 0;
        weight_mem[16'h2F69] <= 0;
        weight_mem[16'h2F6A] <= 0;
        weight_mem[16'h2F6B] <= 0;
        weight_mem[16'h2F6C] <= 0;
        weight_mem[16'h2F6D] <= 0;
        weight_mem[16'h2F6E] <= 0;
        weight_mem[16'h2F6F] <= 0;
        weight_mem[16'h2F70] <= 0;
        weight_mem[16'h2F71] <= 0;
        weight_mem[16'h2F72] <= 0;
        weight_mem[16'h2F73] <= 0;
        weight_mem[16'h2F74] <= 0;
        weight_mem[16'h2F75] <= 0;
        weight_mem[16'h2F76] <= 0;
        weight_mem[16'h2F77] <= 0;
        weight_mem[16'h2F78] <= 0;
        weight_mem[16'h2F79] <= 0;
        weight_mem[16'h2F7A] <= 0;
        weight_mem[16'h2F7B] <= 0;
        weight_mem[16'h2F7C] <= 0;
        weight_mem[16'h2F7D] <= 0;
        weight_mem[16'h2F7E] <= 0;
        weight_mem[16'h2F7F] <= 0;
        weight_mem[16'h2F80] <= 0;
        weight_mem[16'h2F81] <= 0;
        weight_mem[16'h2F82] <= 0;
        weight_mem[16'h2F83] <= 0;
        weight_mem[16'h2F84] <= 0;
        weight_mem[16'h2F85] <= 0;
        weight_mem[16'h2F86] <= 0;
        weight_mem[16'h2F87] <= 0;
        weight_mem[16'h2F88] <= 0;
        weight_mem[16'h2F89] <= 0;
        weight_mem[16'h2F8A] <= 0;
        weight_mem[16'h2F8B] <= 0;
        weight_mem[16'h2F8C] <= 0;
        weight_mem[16'h2F8D] <= 0;
        weight_mem[16'h2F8E] <= 0;
        weight_mem[16'h2F8F] <= 0;
        weight_mem[16'h2F90] <= 0;
        weight_mem[16'h2F91] <= 0;
        weight_mem[16'h2F92] <= 0;
        weight_mem[16'h2F93] <= 0;
        weight_mem[16'h2F94] <= 0;
        weight_mem[16'h2F95] <= 0;
        weight_mem[16'h2F96] <= 0;
        weight_mem[16'h2F97] <= 0;
        weight_mem[16'h2F98] <= 0;
        weight_mem[16'h2F99] <= 0;
        weight_mem[16'h2F9A] <= 0;
        weight_mem[16'h2F9B] <= 0;
        weight_mem[16'h2F9C] <= 0;
        weight_mem[16'h2F9D] <= 0;
        weight_mem[16'h2F9E] <= 0;
        weight_mem[16'h2F9F] <= 0;
        weight_mem[16'h2FA0] <= 0;
        weight_mem[16'h2FA1] <= 0;
        weight_mem[16'h2FA2] <= 0;
        weight_mem[16'h2FA3] <= 0;
        weight_mem[16'h2FA4] <= 0;
        weight_mem[16'h2FA5] <= 0;
        weight_mem[16'h2FA6] <= 0;
        weight_mem[16'h2FA7] <= 0;
        weight_mem[16'h2FA8] <= 0;
        weight_mem[16'h2FA9] <= 0;
        weight_mem[16'h2FAA] <= 0;
        weight_mem[16'h2FAB] <= 0;
        weight_mem[16'h2FAC] <= 0;
        weight_mem[16'h2FAD] <= 0;
        weight_mem[16'h2FAE] <= 0;
        weight_mem[16'h2FAF] <= 0;

        // layer 1 neuron 24
        weight_mem[16'h3000] <= 244;
        weight_mem[16'h3001] <= 4;
        weight_mem[16'h3002] <= 254;
        weight_mem[16'h3003] <= 243;
        weight_mem[16'h3004] <= 255;
        weight_mem[16'h3005] <= 255;
        weight_mem[16'h3006] <= 2;
        weight_mem[16'h3007] <= 246;
        weight_mem[16'h3008] <= 251;
        weight_mem[16'h3009] <= 4;
        weight_mem[16'h300A] <= 2;
        weight_mem[16'h300B] <= 251;
        weight_mem[16'h300C] <= 9;
        weight_mem[16'h300D] <= 247;
        weight_mem[16'h300E] <= 242;
        weight_mem[16'h300F] <= 4;
        weight_mem[16'h3010] <= 6;
        weight_mem[16'h3011] <= 3;
        weight_mem[16'h3012] <= 253;
        weight_mem[16'h3013] <= 7;
        weight_mem[16'h3014] <= 251;
        weight_mem[16'h3015] <= 249;
        weight_mem[16'h3016] <= 242;
        weight_mem[16'h3017] <= 3;
        weight_mem[16'h3018] <= 5;
        weight_mem[16'h3019] <= 2;
        weight_mem[16'h301A] <= 7;
        weight_mem[16'h301B] <= 244;
        weight_mem[16'h301C] <= 250;
        weight_mem[16'h301D] <= 10;
        weight_mem[16'h301E] <= 4;
        weight_mem[16'h301F] <= 243;
        weight_mem[16'h3020] <= 12;
        weight_mem[16'h3021] <= 252;
        weight_mem[16'h3022] <= 12;
        weight_mem[16'h3023] <= 9;
        weight_mem[16'h3024] <= 4;
        weight_mem[16'h3025] <= 14;
        weight_mem[16'h3026] <= 245;
        weight_mem[16'h3027] <= 6;
        weight_mem[16'h3028] <= 251;
        weight_mem[16'h3029] <= 248;
        weight_mem[16'h302A] <= 4;
        weight_mem[16'h302B] <= 8;
        weight_mem[16'h302C] <= 242;
        weight_mem[16'h302D] <= 10;
        weight_mem[16'h302E] <= 1;
        weight_mem[16'h302F] <= 249;
        weight_mem[16'h3030] <= 6;
        weight_mem[16'h3031] <= 253;
        weight_mem[16'h3032] <= 249;
        weight_mem[16'h3033] <= 251;
        weight_mem[16'h3034] <= 248;
        weight_mem[16'h3035] <= 5;
        weight_mem[16'h3036] <= 15;
        weight_mem[16'h3037] <= 21;
        weight_mem[16'h3038] <= 18;
        weight_mem[16'h3039] <= 8;
        weight_mem[16'h303A] <= 13;
        weight_mem[16'h303B] <= 20;
        weight_mem[16'h303C] <= 15;
        weight_mem[16'h303D] <= 15;
        weight_mem[16'h303E] <= 245;
        weight_mem[16'h303F] <= 246;
        weight_mem[16'h3040] <= 9;
        weight_mem[16'h3041] <= 0;
        weight_mem[16'h3042] <= 238;
        weight_mem[16'h3043] <= 237;
        weight_mem[16'h3044] <= 255;
        weight_mem[16'h3045] <= 8;
        weight_mem[16'h3046] <= 8;
        weight_mem[16'h3047] <= 249;
        weight_mem[16'h3048] <= 4;
        weight_mem[16'h3049] <= 5;
        weight_mem[16'h304A] <= 8;
        weight_mem[16'h304B] <= 15;
        weight_mem[16'h304C] <= 18;
        weight_mem[16'h304D] <= 15;
        weight_mem[16'h304E] <= 27;
        weight_mem[16'h304F] <= 18;
        weight_mem[16'h3050] <= 20;
        weight_mem[16'h3051] <= 4;
        weight_mem[16'h3052] <= 13;
        weight_mem[16'h3053] <= 246;
        weight_mem[16'h3054] <= 243;
        weight_mem[16'h3055] <= 245;
        weight_mem[16'h3056] <= 247;
        weight_mem[16'h3057] <= 220;
        weight_mem[16'h3058] <= 223;
        weight_mem[16'h3059] <= 223;
        weight_mem[16'h305A] <= 211;
        weight_mem[16'h305B] <= 214;
        weight_mem[16'h305C] <= 238;
        weight_mem[16'h305D] <= 237;
        weight_mem[16'h305E] <= 4;
        weight_mem[16'h305F] <= 251;
        weight_mem[16'h3060] <= 248;
        weight_mem[16'h3061] <= 247;
        weight_mem[16'h3062] <= 6;
        weight_mem[16'h3063] <= 16;
        weight_mem[16'h3064] <= 15;
        weight_mem[16'h3065] <= 26;
        weight_mem[16'h3066] <= 15;
        weight_mem[16'h3067] <= 241;
        weight_mem[16'h3068] <= 231;
        weight_mem[16'h3069] <= 207;
        weight_mem[16'h306A] <= 202;
        weight_mem[16'h306B] <= 187;
        weight_mem[16'h306C] <= 195;
        weight_mem[16'h306D] <= 219;
        weight_mem[16'h306E] <= 198;
        weight_mem[16'h306F] <= 190;
        weight_mem[16'h3070] <= 196;
        weight_mem[16'h3071] <= 212;
        weight_mem[16'h3072] <= 217;
        weight_mem[16'h3073] <= 207;
        weight_mem[16'h3074] <= 217;
        weight_mem[16'h3075] <= 244;
        weight_mem[16'h3076] <= 1;
        weight_mem[16'h3077] <= 252;
        weight_mem[16'h3078] <= 244;
        weight_mem[16'h3079] <= 9;
        weight_mem[16'h307A] <= 247;
        weight_mem[16'h307B] <= 12;
        weight_mem[16'h307C] <= 25;
        weight_mem[16'h307D] <= 8;
        weight_mem[16'h307E] <= 250;
        weight_mem[16'h307F] <= 244;
        weight_mem[16'h3080] <= 213;
        weight_mem[16'h3081] <= 198;
        weight_mem[16'h3082] <= 182;
        weight_mem[16'h3083] <= 207;
        weight_mem[16'h3084] <= 228;
        weight_mem[16'h3085] <= 242;
        weight_mem[16'h3086] <= 236;
        weight_mem[16'h3087] <= 218;
        weight_mem[16'h3088] <= 244;
        weight_mem[16'h3089] <= 244;
        weight_mem[16'h308A] <= 1;
        weight_mem[16'h308B] <= 241;
        weight_mem[16'h308C] <= 219;
        weight_mem[16'h308D] <= 239;
        weight_mem[16'h308E] <= 244;
        weight_mem[16'h308F] <= 4;
        weight_mem[16'h3090] <= 250;
        weight_mem[16'h3091] <= 6;
        weight_mem[16'h3092] <= 3;
        weight_mem[16'h3093] <= 14;
        weight_mem[16'h3094] <= 19;
        weight_mem[16'h3095] <= 3;
        weight_mem[16'h3096] <= 1;
        weight_mem[16'h3097] <= 212;
        weight_mem[16'h3098] <= 211;
        weight_mem[16'h3099] <= 190;
        weight_mem[16'h309A] <= 175;
        weight_mem[16'h309B] <= 247;
        weight_mem[16'h309C] <= 73;
        weight_mem[16'h309D] <= 91;
        weight_mem[16'h309E] <= 81;
        weight_mem[16'h309F] <= 46;
        weight_mem[16'h30A0] <= 35;
        weight_mem[16'h30A1] <= 52;
        weight_mem[16'h30A2] <= 37;
        weight_mem[16'h30A3] <= 12;
        weight_mem[16'h30A4] <= 246;
        weight_mem[16'h30A5] <= 241;
        weight_mem[16'h30A6] <= 255;
        weight_mem[16'h30A7] <= 5;
        weight_mem[16'h30A8] <= 6;
        weight_mem[16'h30A9] <= 4;
        weight_mem[16'h30AA] <= 4;
        weight_mem[16'h30AB] <= 250;
        weight_mem[16'h30AC] <= 7;
        weight_mem[16'h30AD] <= 241;
        weight_mem[16'h30AE] <= 237;
        weight_mem[16'h30AF] <= 233;
        weight_mem[16'h30B0] <= 231;
        weight_mem[16'h30B1] <= 231;
        weight_mem[16'h30B2] <= 245;
        weight_mem[16'h30B3] <= 38;
        weight_mem[16'h30B4] <= 118;
        weight_mem[16'h30B5] <= 127;
        weight_mem[16'h30B6] <= 82;
        weight_mem[16'h30B7] <= 41;
        weight_mem[16'h30B8] <= 67;
        weight_mem[16'h30B9] <= 86;
        weight_mem[16'h30BA] <= 84;
        weight_mem[16'h30BB] <= 45;
        weight_mem[16'h30BC] <= 248;
        weight_mem[16'h30BD] <= 240;
        weight_mem[16'h30BE] <= 253;
        weight_mem[16'h30BF] <= 250;
        weight_mem[16'h30C0] <= 1;
        weight_mem[16'h30C1] <= 9;
        weight_mem[16'h30C2] <= 243;
        weight_mem[16'h30C3] <= 3;
        weight_mem[16'h30C4] <= 244;
        weight_mem[16'h30C5] <= 248;
        weight_mem[16'h30C6] <= 221;
        weight_mem[16'h30C7] <= 251;
        weight_mem[16'h30C8] <= 245;
        weight_mem[16'h30C9] <= 7;
        weight_mem[16'h30CA] <= 23;
        weight_mem[16'h30CB] <= 46;
        weight_mem[16'h30CC] <= 57;
        weight_mem[16'h30CD] <= 83;
        weight_mem[16'h30CE] <= 51;
        weight_mem[16'h30CF] <= 9;
        weight_mem[16'h30D0] <= 30;
        weight_mem[16'h30D1] <= 71;
        weight_mem[16'h30D2] <= 49;
        weight_mem[16'h30D3] <= 10;
        weight_mem[16'h30D4] <= 232;
        weight_mem[16'h30D5] <= 4;
        weight_mem[16'h30D6] <= 4;
        weight_mem[16'h30D7] <= 2;
        weight_mem[16'h30D8] <= 247;
        weight_mem[16'h30D9] <= 254;
        weight_mem[16'h30DA] <= 3;
        weight_mem[16'h30DB] <= 254;
        weight_mem[16'h30DC] <= 255;
        weight_mem[16'h30DD] <= 241;
        weight_mem[16'h30DE] <= 238;
        weight_mem[16'h30DF] <= 232;
        weight_mem[16'h30E0] <= 235;
        weight_mem[16'h30E1] <= 254;
        weight_mem[16'h30E2] <= 13;
        weight_mem[16'h30E3] <= 45;
        weight_mem[16'h30E4] <= 60;
        weight_mem[16'h30E5] <= 56;
        weight_mem[16'h30E6] <= 54;
        weight_mem[16'h30E7] <= 73;
        weight_mem[16'h30E8] <= 64;
        weight_mem[16'h30E9] <= 42;
        weight_mem[16'h30EA] <= 13;
        weight_mem[16'h30EB] <= 245;
        weight_mem[16'h30EC] <= 230;
        weight_mem[16'h30ED] <= 244;
        weight_mem[16'h30EE] <= 250;
        weight_mem[16'h30EF] <= 8;
        weight_mem[16'h30F0] <= 246;
        weight_mem[16'h30F1] <= 8;
        weight_mem[16'h30F2] <= 6;
        weight_mem[16'h30F3] <= 249;
        weight_mem[16'h30F4] <= 242;
        weight_mem[16'h30F5] <= 0;
        weight_mem[16'h30F6] <= 5;
        weight_mem[16'h30F7] <= 26;
        weight_mem[16'h30F8] <= 9;
        weight_mem[16'h30F9] <= 17;
        weight_mem[16'h30FA] <= 50;
        weight_mem[16'h30FB] <= 70;
        weight_mem[16'h30FC] <= 63;
        weight_mem[16'h30FD] <= 53;
        weight_mem[16'h30FE] <= 52;
        weight_mem[16'h30FF] <= 31;
        weight_mem[16'h3100] <= 25;
        weight_mem[16'h3101] <= 244;
        weight_mem[16'h3102] <= 249;
        weight_mem[16'h3103] <= 233;
        weight_mem[16'h3104] <= 254;
        weight_mem[16'h3105] <= 245;
        weight_mem[16'h3106] <= 246;
        weight_mem[16'h3107] <= 253;
        weight_mem[16'h3108] <= 0;
        weight_mem[16'h3109] <= 245;
        weight_mem[16'h310A] <= 255;
        weight_mem[16'h310B] <= 13;
        weight_mem[16'h310C] <= 3;
        weight_mem[16'h310D] <= 253;
        weight_mem[16'h310E] <= 29;
        weight_mem[16'h310F] <= 52;
        weight_mem[16'h3110] <= 45;
        weight_mem[16'h3111] <= 71;
        weight_mem[16'h3112] <= 92;
        weight_mem[16'h3113] <= 104;
        weight_mem[16'h3114] <= 66;
        weight_mem[16'h3115] <= 40;
        weight_mem[16'h3116] <= 23;
        weight_mem[16'h3117] <= 5;
        weight_mem[16'h3118] <= 245;
        weight_mem[16'h3119] <= 247;
        weight_mem[16'h311A] <= 241;
        weight_mem[16'h311B] <= 239;
        weight_mem[16'h311C] <= 7;
        weight_mem[16'h311D] <= 254;
        weight_mem[16'h311E] <= 245;
        weight_mem[16'h311F] <= 6;
        weight_mem[16'h3120] <= 4;
        weight_mem[16'h3121] <= 2;
        weight_mem[16'h3122] <= 3;
        weight_mem[16'h3123] <= 11;
        weight_mem[16'h3124] <= 251;
        weight_mem[16'h3125] <= 249;
        weight_mem[16'h3126] <= 252;
        weight_mem[16'h3127] <= 17;
        weight_mem[16'h3128] <= 43;
        weight_mem[16'h3129] <= 50;
        weight_mem[16'h312A] <= 64;
        weight_mem[16'h312B] <= 59;
        weight_mem[16'h312C] <= 34;
        weight_mem[16'h312D] <= 24;
        weight_mem[16'h312E] <= 15;
        weight_mem[16'h312F] <= 15;
        weight_mem[16'h3130] <= 8;
        weight_mem[16'h3131] <= 4;
        weight_mem[16'h3132] <= 250;
        weight_mem[16'h3133] <= 245;
        weight_mem[16'h3134] <= 250;
        weight_mem[16'h3135] <= 6;
        weight_mem[16'h3136] <= 248;
        weight_mem[16'h3137] <= 8;
        weight_mem[16'h3138] <= 247;
        weight_mem[16'h3139] <= 245;
        weight_mem[16'h313A] <= 250;
        weight_mem[16'h313B] <= 7;
        weight_mem[16'h313C] <= 2;
        weight_mem[16'h313D] <= 233;
        weight_mem[16'h313E] <= 231;
        weight_mem[16'h313F] <= 222;
        weight_mem[16'h3140] <= 241;
        weight_mem[16'h3141] <= 217;
        weight_mem[16'h3142] <= 205;
        weight_mem[16'h3143] <= 218;
        weight_mem[16'h3144] <= 247;
        weight_mem[16'h3145] <= 236;
        weight_mem[16'h3146] <= 250;
        weight_mem[16'h3147] <= 16;
        weight_mem[16'h3148] <= 4;
        weight_mem[16'h3149] <= 251;
        weight_mem[16'h314A] <= 239;
        weight_mem[16'h314B] <= 240;
        weight_mem[16'h314C] <= 5;
        weight_mem[16'h314D] <= 245;
        weight_mem[16'h314E] <= 247;
        weight_mem[16'h314F] <= 241;
        weight_mem[16'h3150] <= 0;
        weight_mem[16'h3151] <= 246;
        weight_mem[16'h3152] <= 3;
        weight_mem[16'h3153] <= 13;
        weight_mem[16'h3154] <= 7;
        weight_mem[16'h3155] <= 250;
        weight_mem[16'h3156] <= 238;
        weight_mem[16'h3157] <= 223;
        weight_mem[16'h3158] <= 210;
        weight_mem[16'h3159] <= 193;
        weight_mem[16'h315A] <= 192;
        weight_mem[16'h315B] <= 186;
        weight_mem[16'h315C] <= 214;
        weight_mem[16'h315D] <= 211;
        weight_mem[16'h315E] <= 219;
        weight_mem[16'h315F] <= 232;
        weight_mem[16'h3160] <= 235;
        weight_mem[16'h3161] <= 239;
        weight_mem[16'h3162] <= 243;
        weight_mem[16'h3163] <= 236;
        weight_mem[16'h3164] <= 4;
        weight_mem[16'h3165] <= 9;
        weight_mem[16'h3166] <= 249;
        weight_mem[16'h3167] <= 8;
        weight_mem[16'h3168] <= 2;
        weight_mem[16'h3169] <= 247;
        weight_mem[16'h316A] <= 10;
        weight_mem[16'h316B] <= 250;
        weight_mem[16'h316C] <= 253;
        weight_mem[16'h316D] <= 9;
        weight_mem[16'h316E] <= 5;
        weight_mem[16'h316F] <= 0;
        weight_mem[16'h3170] <= 244;
        weight_mem[16'h3171] <= 220;
        weight_mem[16'h3172] <= 229;
        weight_mem[16'h3173] <= 223;
        weight_mem[16'h3174] <= 228;
        weight_mem[16'h3175] <= 245;
        weight_mem[16'h3176] <= 236;
        weight_mem[16'h3177] <= 246;
        weight_mem[16'h3178] <= 247;
        weight_mem[16'h3179] <= 242;
        weight_mem[16'h317A] <= 1;
        weight_mem[16'h317B] <= 248;
        weight_mem[16'h317C] <= 250;
        weight_mem[16'h317D] <= 9;
        weight_mem[16'h317E] <= 6;
        weight_mem[16'h317F] <= 0;
        weight_mem[16'h3180] <= 4;
        weight_mem[16'h3181] <= 248;
        weight_mem[16'h3182] <= 0;
        weight_mem[16'h3183] <= 248;
        weight_mem[16'h3184] <= 244;
        weight_mem[16'h3185] <= 253;
        weight_mem[16'h3186] <= 10;
        weight_mem[16'h3187] <= 254;
        weight_mem[16'h3188] <= 253;
        weight_mem[16'h3189] <= 252;
        weight_mem[16'h318A] <= 10;
        weight_mem[16'h318B] <= 243;
        weight_mem[16'h318C] <= 250;
        weight_mem[16'h318D] <= 2;
        weight_mem[16'h318E] <= 238;
        weight_mem[16'h318F] <= 252;
        weight_mem[16'h3190] <= 244;
        weight_mem[16'h3191] <= 241;
        weight_mem[16'h3192] <= 2;
        weight_mem[16'h3193] <= 242;
        weight_mem[16'h3194] <= 246;
        weight_mem[16'h3195] <= 1;
        weight_mem[16'h3196] <= 3;
        weight_mem[16'h3197] <= 242;
        weight_mem[16'h3198] <= 7;
        weight_mem[16'h3199] <= 2;
        weight_mem[16'h319A] <= 241;
        weight_mem[16'h319B] <= 242;
        weight_mem[16'h319C] <= 252;
        weight_mem[16'h319D] <= 255;
        weight_mem[16'h319E] <= 249;
        weight_mem[16'h319F] <= 255;
        weight_mem[16'h31A0] <= 5;
        weight_mem[16'h31A1] <= 6;
        weight_mem[16'h31A2] <= 244;
        weight_mem[16'h31A3] <= 251;
        weight_mem[16'h31A4] <= 1;
        weight_mem[16'h31A5] <= 245;
        weight_mem[16'h31A6] <= 0;
        weight_mem[16'h31A7] <= 242;
        weight_mem[16'h31A8] <= 5;
        weight_mem[16'h31A9] <= 4;
        weight_mem[16'h31AA] <= 246;
        weight_mem[16'h31AB] <= 0;
        weight_mem[16'h31AC] <= 248;
        weight_mem[16'h31AD] <= 249;
        weight_mem[16'h31AE] <= 10;
        weight_mem[16'h31AF] <= 5;

        // layer 1 neuron 25
        weight_mem[16'h3200] <= 253;
        weight_mem[16'h3201] <= 5;
        weight_mem[16'h3202] <= 243;
        weight_mem[16'h3203] <= 5;
        weight_mem[16'h3204] <= 3;
        weight_mem[16'h3205] <= 250;
        weight_mem[16'h3206] <= 248;
        weight_mem[16'h3207] <= 252;
        weight_mem[16'h3208] <= 254;
        weight_mem[16'h3209] <= 243;
        weight_mem[16'h320A] <= 0;
        weight_mem[16'h320B] <= 252;
        weight_mem[16'h320C] <= 6;
        weight_mem[16'h320D] <= 4;
        weight_mem[16'h320E] <= 5;
        weight_mem[16'h320F] <= 247;
        weight_mem[16'h3210] <= 6;
        weight_mem[16'h3211] <= 6;
        weight_mem[16'h3212] <= 244;
        weight_mem[16'h3213] <= 254;
        weight_mem[16'h3214] <= 4;
        weight_mem[16'h3215] <= 0;
        weight_mem[16'h3216] <= 4;
        weight_mem[16'h3217] <= 243;
        weight_mem[16'h3218] <= 252;
        weight_mem[16'h3219] <= 250;
        weight_mem[16'h321A] <= 253;
        weight_mem[16'h321B] <= 242;
        weight_mem[16'h321C] <= 255;
        weight_mem[16'h321D] <= 7;
        weight_mem[16'h321E] <= 4;
        weight_mem[16'h321F] <= 249;
        weight_mem[16'h3220] <= 2;
        weight_mem[16'h3221] <= 254;
        weight_mem[16'h3222] <= 16;
        weight_mem[16'h3223] <= 12;
        weight_mem[16'h3224] <= 15;
        weight_mem[16'h3225] <= 10;
        weight_mem[16'h3226] <= 253;
        weight_mem[16'h3227] <= 255;
        weight_mem[16'h3228] <= 1;
        weight_mem[16'h3229] <= 252;
        weight_mem[16'h322A] <= 3;
        weight_mem[16'h322B] <= 6;
        weight_mem[16'h322C] <= 6;
        weight_mem[16'h322D] <= 246;
        weight_mem[16'h322E] <= 252;
        weight_mem[16'h322F] <= 243;
        weight_mem[16'h3230] <= 4;
        weight_mem[16'h3231] <= 250;
        weight_mem[16'h3232] <= 5;
        weight_mem[16'h3233] <= 243;
        weight_mem[16'h3234] <= 4;
        weight_mem[16'h3235] <= 253;
        weight_mem[16'h3236] <= 254;
        weight_mem[16'h3237] <= 255;
        weight_mem[16'h3238] <= 18;
        weight_mem[16'h3239] <= 24;
        weight_mem[16'h323A] <= 26;
        weight_mem[16'h323B] <= 30;
        weight_mem[16'h323C] <= 36;
        weight_mem[16'h323D] <= 38;
        weight_mem[16'h323E] <= 27;
        weight_mem[16'h323F] <= 6;
        weight_mem[16'h3240] <= 5;
        weight_mem[16'h3241] <= 1;
        weight_mem[16'h3242] <= 251;
        weight_mem[16'h3243] <= 242;
        weight_mem[16'h3244] <= 2;
        weight_mem[16'h3245] <= 0;
        weight_mem[16'h3246] <= 247;
        weight_mem[16'h3247] <= 255;
        weight_mem[16'h3248] <= 245;
        weight_mem[16'h3249] <= 2;
        weight_mem[16'h324A] <= 247;
        weight_mem[16'h324B] <= 244;
        weight_mem[16'h324C] <= 5;
        weight_mem[16'h324D] <= 11;
        weight_mem[16'h324E] <= 249;
        weight_mem[16'h324F] <= 13;
        weight_mem[16'h3250] <= 255;
        weight_mem[16'h3251] <= 1;
        weight_mem[16'h3252] <= 9;
        weight_mem[16'h3253] <= 29;
        weight_mem[16'h3254] <= 25;
        weight_mem[16'h3255] <= 29;
        weight_mem[16'h3256] <= 23;
        weight_mem[16'h3257] <= 23;
        weight_mem[16'h3258] <= 4;
        weight_mem[16'h3259] <= 246;
        weight_mem[16'h325A] <= 250;
        weight_mem[16'h325B] <= 232;
        weight_mem[16'h325C] <= 238;
        weight_mem[16'h325D] <= 235;
        weight_mem[16'h325E] <= 250;
        weight_mem[16'h325F] <= 5;
        weight_mem[16'h3260] <= 4;
        weight_mem[16'h3261] <= 2;
        weight_mem[16'h3262] <= 244;
        weight_mem[16'h3263] <= 252;
        weight_mem[16'h3264] <= 1;
        weight_mem[16'h3265] <= 255;
        weight_mem[16'h3266] <= 251;
        weight_mem[16'h3267] <= 0;
        weight_mem[16'h3268] <= 247;
        weight_mem[16'h3269] <= 0;
        weight_mem[16'h326A] <= 249;
        weight_mem[16'h326B] <= 231;
        weight_mem[16'h326C] <= 219;
        weight_mem[16'h326D] <= 238;
        weight_mem[16'h326E] <= 246;
        weight_mem[16'h326F] <= 245;
        weight_mem[16'h3270] <= 6;
        weight_mem[16'h3271] <= 252;
        weight_mem[16'h3272] <= 244;
        weight_mem[16'h3273] <= 235;
        weight_mem[16'h3274] <= 231;
        weight_mem[16'h3275] <= 236;
        weight_mem[16'h3276] <= 247;
        weight_mem[16'h3277] <= 6;
        weight_mem[16'h3278] <= 246;
        weight_mem[16'h3279] <= 3;
        weight_mem[16'h327A] <= 6;
        weight_mem[16'h327B] <= 1;
        weight_mem[16'h327C] <= 19;
        weight_mem[16'h327D] <= 10;
        weight_mem[16'h327E] <= 4;
        weight_mem[16'h327F] <= 0;
        weight_mem[16'h3280] <= 15;
        weight_mem[16'h3281] <= 19;
        weight_mem[16'h3282] <= 25;
        weight_mem[16'h3283] <= 44;
        weight_mem[16'h3284] <= 46;
        weight_mem[16'h3285] <= 21;
        weight_mem[16'h3286] <= 237;
        weight_mem[16'h3287] <= 250;
        weight_mem[16'h3288] <= 243;
        weight_mem[16'h3289] <= 240;
        weight_mem[16'h328A] <= 250;
        weight_mem[16'h328B] <= 251;
        weight_mem[16'h328C] <= 244;
        weight_mem[16'h328D] <= 236;
        weight_mem[16'h328E] <= 242;
        weight_mem[16'h328F] <= 251;
        weight_mem[16'h3290] <= 1;
        weight_mem[16'h3291] <= 9;
        weight_mem[16'h3292] <= 10;
        weight_mem[16'h3293] <= 11;
        weight_mem[16'h3294] <= 6;
        weight_mem[16'h3295] <= 7;
        weight_mem[16'h3296] <= 29;
        weight_mem[16'h3297] <= 1;
        weight_mem[16'h3298] <= 4;
        weight_mem[16'h3299] <= 2;
        weight_mem[16'h329A] <= 28;
        weight_mem[16'h329B] <= 93;
        weight_mem[16'h329C] <= 127;
        weight_mem[16'h329D] <= 41;
        weight_mem[16'h329E] <= 16;
        weight_mem[16'h329F] <= 254;
        weight_mem[16'h32A0] <= 252;
        weight_mem[16'h32A1] <= 251;
        weight_mem[16'h32A2] <= 12;
        weight_mem[16'h32A3] <= 8;
        weight_mem[16'h32A4] <= 7;
        weight_mem[16'h32A5] <= 9;
        weight_mem[16'h32A6] <= 7;
        weight_mem[16'h32A7] <= 250;
        weight_mem[16'h32A8] <= 4;
        weight_mem[16'h32A9] <= 3;
        weight_mem[16'h32AA] <= 250;
        weight_mem[16'h32AB] <= 2;
        weight_mem[16'h32AC] <= 8;
        weight_mem[16'h32AD] <= 239;
        weight_mem[16'h32AE] <= 241;
        weight_mem[16'h32AF] <= 212;
        weight_mem[16'h32B0] <= 210;
        weight_mem[16'h32B1] <= 210;
        weight_mem[16'h32B2] <= 3;
        weight_mem[16'h32B3] <= 104;
        weight_mem[16'h32B4] <= 91;
        weight_mem[16'h32B5] <= 7;
        weight_mem[16'h32B6] <= 222;
        weight_mem[16'h32B7] <= 11;
        weight_mem[16'h32B8] <= 22;
        weight_mem[16'h32B9] <= 8;
        weight_mem[16'h32BA] <= 26;
        weight_mem[16'h32BB] <= 24;
        weight_mem[16'h32BC] <= 22;
        weight_mem[16'h32BD] <= 17;
        weight_mem[16'h32BE] <= 8;
        weight_mem[16'h32BF] <= 245;
        weight_mem[16'h32C0] <= 244;
        weight_mem[16'h32C1] <= 0;
        weight_mem[16'h32C2] <= 4;
        weight_mem[16'h32C3] <= 255;
        weight_mem[16'h32C4] <= 236;
        weight_mem[16'h32C5] <= 224;
        weight_mem[16'h32C6] <= 209;
        weight_mem[16'h32C7] <= 201;
        weight_mem[16'h32C8] <= 191;
        weight_mem[16'h32C9] <= 180;
        weight_mem[16'h32CA] <= 227;
        weight_mem[16'h32CB] <= 41;
        weight_mem[16'h32CC] <= 45;
        weight_mem[16'h32CD] <= 230;
        weight_mem[16'h32CE] <= 223;
        weight_mem[16'h32CF] <= 248;
        weight_mem[16'h32D0] <= 248;
        weight_mem[16'h32D1] <= 245;
        weight_mem[16'h32D2] <= 2;
        weight_mem[16'h32D3] <= 24;
        weight_mem[16'h32D4] <= 32;
        weight_mem[16'h32D5] <= 3;
        weight_mem[16'h32D6] <= 249;
        weight_mem[16'h32D7] <= 5;
        weight_mem[16'h32D8] <= 246;
        weight_mem[16'h32D9] <= 248;
        weight_mem[16'h32DA] <= 0;
        weight_mem[16'h32DB] <= 249;
        weight_mem[16'h32DC] <= 219;
        weight_mem[16'h32DD] <= 201;
        weight_mem[16'h32DE] <= 197;
        weight_mem[16'h32DF] <= 183;
        weight_mem[16'h32E0] <= 199;
        weight_mem[16'h32E1] <= 177;
        weight_mem[16'h32E2] <= 193;
        weight_mem[16'h32E3] <= 8;
        weight_mem[16'h32E4] <= 24;
        weight_mem[16'h32E5] <= 3;
        weight_mem[16'h32E6] <= 221;
        weight_mem[16'h32E7] <= 229;
        weight_mem[16'h32E8] <= 248;
        weight_mem[16'h32E9] <= 254;
        weight_mem[16'h32EA] <= 14;
        weight_mem[16'h32EB] <= 6;
        weight_mem[16'h32EC] <= 15;
        weight_mem[16'h32ED] <= 7;
        weight_mem[16'h32EE] <= 249;
        weight_mem[16'h32EF] <= 254;
        weight_mem[16'h32F0] <= 245;
        weight_mem[16'h32F1] <= 2;
        weight_mem[16'h32F2] <= 2;
        weight_mem[16'h32F3] <= 253;
        weight_mem[16'h32F4] <= 248;
        weight_mem[16'h32F5] <= 234;
        weight_mem[16'h32F6] <= 208;
        weight_mem[16'h32F7] <= 196;
        weight_mem[16'h32F8] <= 205;
        weight_mem[16'h32F9] <= 212;
        weight_mem[16'h32FA] <= 207;
        weight_mem[16'h32FB] <= 245;
        weight_mem[16'h32FC] <= 20;
        weight_mem[16'h32FD] <= 209;
        weight_mem[16'h32FE] <= 182;
        weight_mem[16'h32FF] <= 199;
        weight_mem[16'h3300] <= 244;
        weight_mem[16'h3301] <= 3;
        weight_mem[16'h3302] <= 18;
        weight_mem[16'h3303] <= 9;
        weight_mem[16'h3304] <= 21;
        weight_mem[16'h3305] <= 27;
        weight_mem[16'h3306] <= 10;
        weight_mem[16'h3307] <= 249;
        weight_mem[16'h3308] <= 5;
        weight_mem[16'h3309] <= 2;
        weight_mem[16'h330A] <= 248;
        weight_mem[16'h330B] <= 253;
        weight_mem[16'h330C] <= 17;
        weight_mem[16'h330D] <= 249;
        weight_mem[16'h330E] <= 7;
        weight_mem[16'h330F] <= 8;
        weight_mem[16'h3310] <= 5;
        weight_mem[16'h3311] <= 16;
        weight_mem[16'h3312] <= 246;
        weight_mem[16'h3313] <= 239;
        weight_mem[16'h3314] <= 245;
        weight_mem[16'h3315] <= 207;
        weight_mem[16'h3316] <= 206;
        weight_mem[16'h3317] <= 241;
        weight_mem[16'h3318] <= 255;
        weight_mem[16'h3319] <= 24;
        weight_mem[16'h331A] <= 24;
        weight_mem[16'h331B] <= 41;
        weight_mem[16'h331C] <= 17;
        weight_mem[16'h331D] <= 21;
        weight_mem[16'h331E] <= 249;
        weight_mem[16'h331F] <= 247;
        weight_mem[16'h3320] <= 254;
        weight_mem[16'h3321] <= 244;
        weight_mem[16'h3322] <= 254;
        weight_mem[16'h3323] <= 18;
        weight_mem[16'h3324] <= 26;
        weight_mem[16'h3325] <= 18;
        weight_mem[16'h3326] <= 45;
        weight_mem[16'h3327] <= 72;
        weight_mem[16'h3328] <= 71;
        weight_mem[16'h3329] <= 71;
        weight_mem[16'h332A] <= 69;
        weight_mem[16'h332B] <= 56;
        weight_mem[16'h332C] <= 19;
        weight_mem[16'h332D] <= 252;
        weight_mem[16'h332E] <= 254;
        weight_mem[16'h332F] <= 2;
        weight_mem[16'h3330] <= 12;
        weight_mem[16'h3331] <= 9;
        weight_mem[16'h3332] <= 21;
        weight_mem[16'h3333] <= 31;
        weight_mem[16'h3334] <= 21;
        weight_mem[16'h3335] <= 15;
        weight_mem[16'h3336] <= 9;
        weight_mem[16'h3337] <= 243;
        weight_mem[16'h3338] <= 4;
        weight_mem[16'h3339] <= 243;
        weight_mem[16'h333A] <= 254;
        weight_mem[16'h333B] <= 18;
        weight_mem[16'h333C] <= 30;
        weight_mem[16'h333D] <= 34;
        weight_mem[16'h333E] <= 50;
        weight_mem[16'h333F] <= 69;
        weight_mem[16'h3340] <= 63;
        weight_mem[16'h3341] <= 69;
        weight_mem[16'h3342] <= 74;
        weight_mem[16'h3343] <= 43;
        weight_mem[16'h3344] <= 41;
        weight_mem[16'h3345] <= 2;
        weight_mem[16'h3346] <= 251;
        weight_mem[16'h3347] <= 248;
        weight_mem[16'h3348] <= 1;
        weight_mem[16'h3349] <= 253;
        weight_mem[16'h334A] <= 254;
        weight_mem[16'h334B] <= 251;
        weight_mem[16'h334C] <= 3;
        weight_mem[16'h334D] <= 250;
        weight_mem[16'h334E] <= 243;
        weight_mem[16'h334F] <= 254;
        weight_mem[16'h3350] <= 5;
        weight_mem[16'h3351] <= 3;
        weight_mem[16'h3352] <= 9;
        weight_mem[16'h3353] <= 255;
        weight_mem[16'h3354] <= 20;
        weight_mem[16'h3355] <= 34;
        weight_mem[16'h3356] <= 36;
        weight_mem[16'h3357] <= 30;
        weight_mem[16'h3358] <= 24;
        weight_mem[16'h3359] <= 22;
        weight_mem[16'h335A] <= 25;
        weight_mem[16'h335B] <= 35;
        weight_mem[16'h335C] <= 15;
        weight_mem[16'h335D] <= 3;
        weight_mem[16'h335E] <= 239;
        weight_mem[16'h335F] <= 225;
        weight_mem[16'h3360] <= 231;
        weight_mem[16'h3361] <= 235;
        weight_mem[16'h3362] <= 237;
        weight_mem[16'h3363] <= 254;
        weight_mem[16'h3364] <= 243;
        weight_mem[16'h3365] <= 247;
        weight_mem[16'h3366] <= 0;
        weight_mem[16'h3367] <= 1;
        weight_mem[16'h3368] <= 2;
        weight_mem[16'h3369] <= 7;
        weight_mem[16'h336A] <= 244;
        weight_mem[16'h336B] <= 254;
        weight_mem[16'h336C] <= 250;
        weight_mem[16'h336D] <= 11;
        weight_mem[16'h336E] <= 255;
        weight_mem[16'h336F] <= 15;
        weight_mem[16'h3370] <= 254;
        weight_mem[16'h3371] <= 241;
        weight_mem[16'h3372] <= 254;
        weight_mem[16'h3373] <= 11;
        weight_mem[16'h3374] <= 14;
        weight_mem[16'h3375] <= 7;
        weight_mem[16'h3376] <= 245;
        weight_mem[16'h3377] <= 239;
        weight_mem[16'h3378] <= 242;
        weight_mem[16'h3379] <= 245;
        weight_mem[16'h337A] <= 235;
        weight_mem[16'h337B] <= 0;
        weight_mem[16'h337C] <= 240;
        weight_mem[16'h337D] <= 253;
        weight_mem[16'h337E] <= 246;
        weight_mem[16'h337F] <= 243;
        weight_mem[16'h3380] <= 249;
        weight_mem[16'h3381] <= 244;
        weight_mem[16'h3382] <= 253;
        weight_mem[16'h3383] <= 246;
        weight_mem[16'h3384] <= 250;
        weight_mem[16'h3385] <= 5;
        weight_mem[16'h3386] <= 1;
        weight_mem[16'h3387] <= 250;
        weight_mem[16'h3388] <= 247;
        weight_mem[16'h3389] <= 5;
        weight_mem[16'h338A] <= 9;
        weight_mem[16'h338B] <= 5;
        weight_mem[16'h338C] <= 16;
        weight_mem[16'h338D] <= 16;
        weight_mem[16'h338E] <= 18;
        weight_mem[16'h338F] <= 14;
        weight_mem[16'h3390] <= 243;
        weight_mem[16'h3391] <= 242;
        weight_mem[16'h3392] <= 247;
        weight_mem[16'h3393] <= 4;
        weight_mem[16'h3394] <= 253;
        weight_mem[16'h3395] <= 1;
        weight_mem[16'h3396] <= 254;
        weight_mem[16'h3397] <= 255;
        weight_mem[16'h3398] <= 3;
        weight_mem[16'h3399] <= 4;
        weight_mem[16'h339A] <= 0;
        weight_mem[16'h339B] <= 241;
        weight_mem[16'h339C] <= 254;
        weight_mem[16'h339D] <= 253;
        weight_mem[16'h339E] <= 245;
        weight_mem[16'h339F] <= 6;
        weight_mem[16'h33A0] <= 255;
        weight_mem[16'h33A1] <= 251;
        weight_mem[16'h33A2] <= 249;
        weight_mem[16'h33A3] <= 6;
        weight_mem[16'h33A4] <= 254;
        weight_mem[16'h33A5] <= 249;
        weight_mem[16'h33A6] <= 3;
        weight_mem[16'h33A7] <= 8;
        weight_mem[16'h33A8] <= 1;
        weight_mem[16'h33A9] <= 3;
        weight_mem[16'h33AA] <= 252;
        weight_mem[16'h33AB] <= 246;
        weight_mem[16'h33AC] <= 246;
        weight_mem[16'h33AD] <= 243;
        weight_mem[16'h33AE] <= 3;
        weight_mem[16'h33AF] <= 253;

        // layer 1 neuron 26
        weight_mem[16'h3400] <= 249;
        weight_mem[16'h3401] <= 3;
        weight_mem[16'h3402] <= 247;
        weight_mem[16'h3403] <= 246;
        weight_mem[16'h3404] <= 0;
        weight_mem[16'h3405] <= 247;
        weight_mem[16'h3406] <= 3;
        weight_mem[16'h3407] <= 3;
        weight_mem[16'h3408] <= 8;
        weight_mem[16'h3409] <= 4;
        weight_mem[16'h340A] <= 251;
        weight_mem[16'h340B] <= 255;
        weight_mem[16'h340C] <= 2;
        weight_mem[16'h340D] <= 250;
        weight_mem[16'h340E] <= 4;
        weight_mem[16'h340F] <= 1;
        weight_mem[16'h3410] <= 2;
        weight_mem[16'h3411] <= 1;
        weight_mem[16'h3412] <= 252;
        weight_mem[16'h3413] <= 0;
        weight_mem[16'h3414] <= 1;
        weight_mem[16'h3415] <= 248;
        weight_mem[16'h3416] <= 3;
        weight_mem[16'h3417] <= 8;
        weight_mem[16'h3418] <= 246;
        weight_mem[16'h3419] <= 248;
        weight_mem[16'h341A] <= 6;
        weight_mem[16'h341B] <= 7;
        weight_mem[16'h341C] <= 251;
        weight_mem[16'h341D] <= 9;
        weight_mem[16'h341E] <= 248;
        weight_mem[16'h341F] <= 248;
        weight_mem[16'h3420] <= 246;
        weight_mem[16'h3421] <= 5;
        weight_mem[16'h3422] <= 249;
        weight_mem[16'h3423] <= 250;
        weight_mem[16'h3424] <= 247;
        weight_mem[16'h3425] <= 242;
        weight_mem[16'h3426] <= 1;
        weight_mem[16'h3427] <= 255;
        weight_mem[16'h3428] <= 255;
        weight_mem[16'h3429] <= 1;
        weight_mem[16'h342A] <= 251;
        weight_mem[16'h342B] <= 251;
        weight_mem[16'h342C] <= 252;
        weight_mem[16'h342D] <= 251;
        weight_mem[16'h342E] <= 6;
        weight_mem[16'h342F] <= 246;
        weight_mem[16'h3430] <= 6;
        weight_mem[16'h3431] <= 255;
        weight_mem[16'h3432] <= 248;
        weight_mem[16'h3433] <= 251;
        weight_mem[16'h3434] <= 252;
        weight_mem[16'h3435] <= 248;
        weight_mem[16'h3436] <= 6;
        weight_mem[16'h3437] <= 3;
        weight_mem[16'h3438] <= 254;
        weight_mem[16'h3439] <= 241;
        weight_mem[16'h343A] <= 236;
        weight_mem[16'h343B] <= 227;
        weight_mem[16'h343C] <= 240;
        weight_mem[16'h343D] <= 227;
        weight_mem[16'h343E] <= 227;
        weight_mem[16'h343F] <= 243;
        weight_mem[16'h3440] <= 245;
        weight_mem[16'h3441] <= 252;
        weight_mem[16'h3442] <= 255;
        weight_mem[16'h3443] <= 1;
        weight_mem[16'h3444] <= 0;
        weight_mem[16'h3445] <= 251;
        weight_mem[16'h3446] <= 254;
        weight_mem[16'h3447] <= 5;
        weight_mem[16'h3448] <= 249;
        weight_mem[16'h3449] <= 6;
        weight_mem[16'h344A] <= 7;
        weight_mem[16'h344B] <= 1;
        weight_mem[16'h344C] <= 248;
        weight_mem[16'h344D] <= 249;
        weight_mem[16'h344E] <= 1;
        weight_mem[16'h344F] <= 249;
        weight_mem[16'h3450] <= 240;
        weight_mem[16'h3451] <= 4;
        weight_mem[16'h3452] <= 252;
        weight_mem[16'h3453] <= 12;
        weight_mem[16'h3454] <= 244;
        weight_mem[16'h3455] <= 238;
        weight_mem[16'h3456] <= 0;
        weight_mem[16'h3457] <= 3;
        weight_mem[16'h3458] <= 238;
        weight_mem[16'h3459] <= 248;
        weight_mem[16'h345A] <= 255;
        weight_mem[16'h345B] <= 252;
        weight_mem[16'h345C] <= 3;
        weight_mem[16'h345D] <= 10;
        weight_mem[16'h345E] <= 247;
        weight_mem[16'h345F] <= 2;
        weight_mem[16'h3460] <= 3;
        weight_mem[16'h3461] <= 249;
        weight_mem[16'h3462] <= 4;
        weight_mem[16'h3463] <= 254;
        weight_mem[16'h3464] <= 241;
        weight_mem[16'h3465] <= 253;
        weight_mem[16'h3466] <= 253;
        weight_mem[16'h3467] <= 252;
        weight_mem[16'h3468] <= 240;
        weight_mem[16'h3469] <= 244;
        weight_mem[16'h346A] <= 236;
        weight_mem[16'h346B] <= 228;
        weight_mem[16'h346C] <= 239;
        weight_mem[16'h346D] <= 244;
        weight_mem[16'h346E] <= 229;
        weight_mem[16'h346F] <= 225;
        weight_mem[16'h3470] <= 234;
        weight_mem[16'h3471] <= 239;
        weight_mem[16'h3472] <= 238;
        weight_mem[16'h3473] <= 1;
        weight_mem[16'h3474] <= 16;
        weight_mem[16'h3475] <= 6;
        weight_mem[16'h3476] <= 0;
        weight_mem[16'h3477] <= 5;
        weight_mem[16'h3478] <= 1;
        weight_mem[16'h3479] <= 1;
        weight_mem[16'h347A] <= 3;
        weight_mem[16'h347B] <= 247;
        weight_mem[16'h347C] <= 246;
        weight_mem[16'h347D] <= 242;
        weight_mem[16'h347E] <= 245;
        weight_mem[16'h347F] <= 236;
        weight_mem[16'h3480] <= 229;
        weight_mem[16'h3481] <= 218;
        weight_mem[16'h3482] <= 226;
        weight_mem[16'h3483] <= 251;
        weight_mem[16'h3484] <= 252;
        weight_mem[16'h3485] <= 234;
        weight_mem[16'h3486] <= 210;
        weight_mem[16'h3487] <= 219;
        weight_mem[16'h3488] <= 216;
        weight_mem[16'h3489] <= 243;
        weight_mem[16'h348A] <= 249;
        weight_mem[16'h348B] <= 13;
        weight_mem[16'h348C] <= 28;
        weight_mem[16'h348D] <= 28;
        weight_mem[16'h348E] <= 254;
        weight_mem[16'h348F] <= 8;
        weight_mem[16'h3490] <= 252;
        weight_mem[16'h3491] <= 253;
        weight_mem[16'h3492] <= 254;
        weight_mem[16'h3493] <= 3;
        weight_mem[16'h3494] <= 16;
        weight_mem[16'h3495] <= 8;
        weight_mem[16'h3496] <= 19;
        weight_mem[16'h3497] <= 11;
        weight_mem[16'h3498] <= 9;
        weight_mem[16'h3499] <= 37;
        weight_mem[16'h349A] <= 76;
        weight_mem[16'h349B] <= 124;
        weight_mem[16'h349C] <= 79;
        weight_mem[16'h349D] <= 233;
        weight_mem[16'h349E] <= 203;
        weight_mem[16'h349F] <= 227;
        weight_mem[16'h34A0] <= 250;
        weight_mem[16'h34A1] <= 10;
        weight_mem[16'h34A2] <= 3;
        weight_mem[16'h34A3] <= 22;
        weight_mem[16'h34A4] <= 25;
        weight_mem[16'h34A5] <= 5;
        weight_mem[16'h34A6] <= 249;
        weight_mem[16'h34A7] <= 253;
        weight_mem[16'h34A8] <= 7;
        weight_mem[16'h34A9] <= 255;
        weight_mem[16'h34AA] <= 246;
        weight_mem[16'h34AB] <= 2;
        weight_mem[16'h34AC] <= 36;
        weight_mem[16'h34AD] <= 52;
        weight_mem[16'h34AE] <= 61;
        weight_mem[16'h34AF] <= 70;
        weight_mem[16'h34B0] <= 91;
        weight_mem[16'h34B1] <= 97;
        weight_mem[16'h34B2] <= 115;
        weight_mem[16'h34B3] <= 127;
        weight_mem[16'h34B4] <= 64;
        weight_mem[16'h34B5] <= 230;
        weight_mem[16'h34B6] <= 228;
        weight_mem[16'h34B7] <= 255;
        weight_mem[16'h34B8] <= 3;
        weight_mem[16'h34B9] <= 2;
        weight_mem[16'h34BA] <= 15;
        weight_mem[16'h34BB] <= 15;
        weight_mem[16'h34BC] <= 14;
        weight_mem[16'h34BD] <= 11;
        weight_mem[16'h34BE] <= 250;
        weight_mem[16'h34BF] <= 254;
        weight_mem[16'h34C0] <= 253;
        weight_mem[16'h34C1] <= 0;
        weight_mem[16'h34C2] <= 4;
        weight_mem[16'h34C3] <= 15;
        weight_mem[16'h34C4] <= 40;
        weight_mem[16'h34C5] <= 62;
        weight_mem[16'h34C6] <= 85;
        weight_mem[16'h34C7] <= 81;
        weight_mem[16'h34C8] <= 65;
        weight_mem[16'h34C9] <= 47;
        weight_mem[16'h34CA] <= 33;
        weight_mem[16'h34CB] <= 21;
        weight_mem[16'h34CC] <= 254;
        weight_mem[16'h34CD] <= 236;
        weight_mem[16'h34CE] <= 251;
        weight_mem[16'h34CF] <= 0;
        weight_mem[16'h34D0] <= 24;
        weight_mem[16'h34D1] <= 24;
        weight_mem[16'h34D2] <= 7;
        weight_mem[16'h34D3] <= 20;
        weight_mem[16'h34D4] <= 6;
        weight_mem[16'h34D5] <= 254;
        weight_mem[16'h34D6] <= 246;
        weight_mem[16'h34D7] <= 248;
        weight_mem[16'h34D8] <= 9;
        weight_mem[16'h34D9] <= 1;
        weight_mem[16'h34DA] <= 250;
        weight_mem[16'h34DB] <= 254;
        weight_mem[16'h34DC] <= 34;
        weight_mem[16'h34DD] <= 46;
        weight_mem[16'h34DE] <= 24;
        weight_mem[16'h34DF] <= 15;
        weight_mem[16'h34E0] <= 246;
        weight_mem[16'h34E1] <= 232;
        weight_mem[16'h34E2] <= 227;
        weight_mem[16'h34E3] <= 224;
        weight_mem[16'h34E4] <= 213;
        weight_mem[16'h34E5] <= 231;
        weight_mem[16'h34E6] <= 248;
        weight_mem[16'h34E7] <= 5;
        weight_mem[16'h34E8] <= 7;
        weight_mem[16'h34E9] <= 254;
        weight_mem[16'h34EA] <= 5;
        weight_mem[16'h34EB] <= 9;
        weight_mem[16'h34EC] <= 3;
        weight_mem[16'h34ED] <= 252;
        weight_mem[16'h34EE] <= 5;
        weight_mem[16'h34EF] <= 255;
        weight_mem[16'h34F0] <= 7;
        weight_mem[16'h34F1] <= 4;
        weight_mem[16'h34F2] <= 254;
        weight_mem[16'h34F3] <= 243;
        weight_mem[16'h34F4] <= 249;
        weight_mem[16'h34F5] <= 250;
        weight_mem[16'h34F6] <= 233;
        weight_mem[16'h34F7] <= 244;
        weight_mem[16'h34F8] <= 224;
        weight_mem[16'h34F9] <= 233;
        weight_mem[16'h34FA] <= 232;
        weight_mem[16'h34FB] <= 217;
        weight_mem[16'h34FC] <= 225;
        weight_mem[16'h34FD] <= 0;
        weight_mem[16'h34FE] <= 19;
        weight_mem[16'h34FF] <= 251;
        weight_mem[16'h3500] <= 243;
        weight_mem[16'h3501] <= 2;
        weight_mem[16'h3502] <= 2;
        weight_mem[16'h3503] <= 11;
        weight_mem[16'h3504] <= 252;
        weight_mem[16'h3505] <= 245;
        weight_mem[16'h3506] <= 248;
        weight_mem[16'h3507] <= 3;
        weight_mem[16'h3508] <= 7;
        weight_mem[16'h3509] <= 250;
        weight_mem[16'h350A] <= 3;
        weight_mem[16'h350B] <= 242;
        weight_mem[16'h350C] <= 231;
        weight_mem[16'h350D] <= 242;
        weight_mem[16'h350E] <= 245;
        weight_mem[16'h350F] <= 247;
        weight_mem[16'h3510] <= 247;
        weight_mem[16'h3511] <= 3;
        weight_mem[16'h3512] <= 239;
        weight_mem[16'h3513] <= 218;
        weight_mem[16'h3514] <= 2;
        weight_mem[16'h3515] <= 22;
        weight_mem[16'h3516] <= 14;
        weight_mem[16'h3517] <= 253;
        weight_mem[16'h3518] <= 4;
        weight_mem[16'h3519] <= 6;
        weight_mem[16'h351A] <= 7;
        weight_mem[16'h351B] <= 250;
        weight_mem[16'h351C] <= 247;
        weight_mem[16'h351D] <= 239;
        weight_mem[16'h351E] <= 4;
        weight_mem[16'h351F] <= 5;
        weight_mem[16'h3520] <= 255;
        weight_mem[16'h3521] <= 251;
        weight_mem[16'h3522] <= 251;
        weight_mem[16'h3523] <= 235;
        weight_mem[16'h3524] <= 238;
        weight_mem[16'h3525] <= 249;
        weight_mem[16'h3526] <= 254;
        weight_mem[16'h3527] <= 249;
        weight_mem[16'h3528] <= 6;
        weight_mem[16'h3529] <= 252;
        weight_mem[16'h352A] <= 244;
        weight_mem[16'h352B] <= 243;
        weight_mem[16'h352C] <= 19;
        weight_mem[16'h352D] <= 20;
        weight_mem[16'h352E] <= 252;
        weight_mem[16'h352F] <= 249;
        weight_mem[16'h3530] <= 246;
        weight_mem[16'h3531] <= 4;
        weight_mem[16'h3532] <= 249;
        weight_mem[16'h3533] <= 247;
        weight_mem[16'h3534] <= 247;
        weight_mem[16'h3535] <= 240;
        weight_mem[16'h3536] <= 248;
        weight_mem[16'h3537] <= 2;
        weight_mem[16'h3538] <= 250;
        weight_mem[16'h3539] <= 250;
        weight_mem[16'h353A] <= 254;
        weight_mem[16'h353B] <= 227;
        weight_mem[16'h353C] <= 229;
        weight_mem[16'h353D] <= 238;
        weight_mem[16'h353E] <= 248;
        weight_mem[16'h353F] <= 243;
        weight_mem[16'h3540] <= 248;
        weight_mem[16'h3541] <= 252;
        weight_mem[16'h3542] <= 5;
        weight_mem[16'h3543] <= 11;
        weight_mem[16'h3544] <= 2;
        weight_mem[16'h3545] <= 5;
        weight_mem[16'h3546] <= 5;
        weight_mem[16'h3547] <= 2;
        weight_mem[16'h3548] <= 254;
        weight_mem[16'h3549] <= 248;
        weight_mem[16'h354A] <= 255;
        weight_mem[16'h354B] <= 242;
        weight_mem[16'h354C] <= 239;
        weight_mem[16'h354D] <= 252;
        weight_mem[16'h354E] <= 6;
        weight_mem[16'h354F] <= 5;
        weight_mem[16'h3550] <= 254;
        weight_mem[16'h3551] <= 246;
        weight_mem[16'h3552] <= 250;
        weight_mem[16'h3553] <= 249;
        weight_mem[16'h3554] <= 235;
        weight_mem[16'h3555] <= 226;
        weight_mem[16'h3556] <= 237;
        weight_mem[16'h3557] <= 11;
        weight_mem[16'h3558] <= 0;
        weight_mem[16'h3559] <= 9;
        weight_mem[16'h355A] <= 26;
        weight_mem[16'h355B] <= 13;
        weight_mem[16'h355C] <= 4;
        weight_mem[16'h355D] <= 255;
        weight_mem[16'h355E] <= 8;
        weight_mem[16'h355F] <= 250;
        weight_mem[16'h3560] <= 254;
        weight_mem[16'h3561] <= 6;
        weight_mem[16'h3562] <= 253;
        weight_mem[16'h3563] <= 251;
        weight_mem[16'h3564] <= 248;
        weight_mem[16'h3565] <= 4;
        weight_mem[16'h3566] <= 255;
        weight_mem[16'h3567] <= 9;
        weight_mem[16'h3568] <= 250;
        weight_mem[16'h3569] <= 252;
        weight_mem[16'h356A] <= 250;
        weight_mem[16'h356B] <= 243;
        weight_mem[16'h356C] <= 232;
        weight_mem[16'h356D] <= 226;
        weight_mem[16'h356E] <= 242;
        weight_mem[16'h356F] <= 1;
        weight_mem[16'h3570] <= 255;
        weight_mem[16'h3571] <= 255;
        weight_mem[16'h3572] <= 1;
        weight_mem[16'h3573] <= 245;
        weight_mem[16'h3574] <= 9;
        weight_mem[16'h3575] <= 1;
        weight_mem[16'h3576] <= 17;
        weight_mem[16'h3577] <= 11;
        weight_mem[16'h3578] <= 17;
        weight_mem[16'h3579] <= 16;
        weight_mem[16'h357A] <= 16;
        weight_mem[16'h357B] <= 11;
        weight_mem[16'h357C] <= 251;
        weight_mem[16'h357D] <= 245;
        weight_mem[16'h357E] <= 4;
        weight_mem[16'h357F] <= 246;
        weight_mem[16'h3580] <= 0;
        weight_mem[16'h3581] <= 4;
        weight_mem[16'h3582] <= 1;
        weight_mem[16'h3583] <= 248;
        weight_mem[16'h3584] <= 246;
        weight_mem[16'h3585] <= 250;
        weight_mem[16'h3586] <= 1;
        weight_mem[16'h3587] <= 250;
        weight_mem[16'h3588] <= 239;
        weight_mem[16'h3589] <= 238;
        weight_mem[16'h358A] <= 227;
        weight_mem[16'h358B] <= 227;
        weight_mem[16'h358C] <= 251;
        weight_mem[16'h358D] <= 255;
        weight_mem[16'h358E] <= 252;
        weight_mem[16'h358F] <= 2;
        weight_mem[16'h3590] <= 16;
        weight_mem[16'h3591] <= 8;
        weight_mem[16'h3592] <= 1;
        weight_mem[16'h3593] <= 2;
        weight_mem[16'h3594] <= 9;
        weight_mem[16'h3595] <= 252;
        weight_mem[16'h3596] <= 250;
        weight_mem[16'h3597] <= 255;
        weight_mem[16'h3598] <= 246;
        weight_mem[16'h3599] <= 254;
        weight_mem[16'h359A] <= 255;
        weight_mem[16'h359B] <= 2;
        weight_mem[16'h359C] <= 248;
        weight_mem[16'h359D] <= 249;
        weight_mem[16'h359E] <= 5;
        weight_mem[16'h359F] <= 8;
        weight_mem[16'h35A0] <= 245;
        weight_mem[16'h35A1] <= 1;
        weight_mem[16'h35A2] <= 253;
        weight_mem[16'h35A3] <= 248;
        weight_mem[16'h35A4] <= 245;
        weight_mem[16'h35A5] <= 1;
        weight_mem[16'h35A6] <= 252;
        weight_mem[16'h35A7] <= 252;
        weight_mem[16'h35A8] <= 0;
        weight_mem[16'h35A9] <= 251;
        weight_mem[16'h35AA] <= 255;
        weight_mem[16'h35AB] <= 2;
        weight_mem[16'h35AC] <= 250;
        weight_mem[16'h35AD] <= 4;
        weight_mem[16'h35AE] <= 251;
        weight_mem[16'h35AF] <= 6;

        // layer 1 neuron 27
        weight_mem[16'h3600] <= 0;
        weight_mem[16'h3601] <= 4;
        weight_mem[16'h3602] <= 7;
        weight_mem[16'h3603] <= 255;
        weight_mem[16'h3604] <= 253;
        weight_mem[16'h3605] <= 6;
        weight_mem[16'h3606] <= 1;
        weight_mem[16'h3607] <= 252;
        weight_mem[16'h3608] <= 255;
        weight_mem[16'h3609] <= 251;
        weight_mem[16'h360A] <= 0;
        weight_mem[16'h360B] <= 9;
        weight_mem[16'h360C] <= 254;
        weight_mem[16'h360D] <= 251;
        weight_mem[16'h360E] <= 255;
        weight_mem[16'h360F] <= 253;
        weight_mem[16'h3610] <= 7;
        weight_mem[16'h3611] <= 9;
        weight_mem[16'h3612] <= 12;
        weight_mem[16'h3613] <= 255;
        weight_mem[16'h3614] <= 248;
        weight_mem[16'h3615] <= 5;
        weight_mem[16'h3616] <= 3;
        weight_mem[16'h3617] <= 8;
        weight_mem[16'h3618] <= 0;
        weight_mem[16'h3619] <= 253;
        weight_mem[16'h361A] <= 10;
        weight_mem[16'h361B] <= 10;
        weight_mem[16'h361C] <= 252;
        weight_mem[16'h361D] <= 12;
        weight_mem[16'h361E] <= 11;
        weight_mem[16'h361F] <= 3;
        weight_mem[16'h3620] <= 3;
        weight_mem[16'h3621] <= 247;
        weight_mem[16'h3622] <= 241;
        weight_mem[16'h3623] <= 243;
        weight_mem[16'h3624] <= 246;
        weight_mem[16'h3625] <= 6;
        weight_mem[16'h3626] <= 255;
        weight_mem[16'h3627] <= 4;
        weight_mem[16'h3628] <= 247;
        weight_mem[16'h3629] <= 253;
        weight_mem[16'h362A] <= 252;
        weight_mem[16'h362B] <= 10;
        weight_mem[16'h362C] <= 1;
        weight_mem[16'h362D] <= 8;
        weight_mem[16'h362E] <= 10;
        weight_mem[16'h362F] <= 251;
        weight_mem[16'h3630] <= 250;
        weight_mem[16'h3631] <= 0;
        weight_mem[16'h3632] <= 251;
        weight_mem[16'h3633] <= 251;
        weight_mem[16'h3634] <= 255;
        weight_mem[16'h3635] <= 255;
        weight_mem[16'h3636] <= 7;
        weight_mem[16'h3637] <= 3;
        weight_mem[16'h3638] <= 2;
        weight_mem[16'h3639] <= 5;
        weight_mem[16'h363A] <= 249;
        weight_mem[16'h363B] <= 4;
        weight_mem[16'h363C] <= 6;
        weight_mem[16'h363D] <= 7;
        weight_mem[16'h363E] <= 3;
        weight_mem[16'h363F] <= 5;
        weight_mem[16'h3640] <= 249;
        weight_mem[16'h3641] <= 17;
        weight_mem[16'h3642] <= 5;
        weight_mem[16'h3643] <= 9;
        weight_mem[16'h3644] <= 0;
        weight_mem[16'h3645] <= 12;
        weight_mem[16'h3646] <= 249;
        weight_mem[16'h3647] <= 255;
        weight_mem[16'h3648] <= 250;
        weight_mem[16'h3649] <= 10;
        weight_mem[16'h364A] <= 252;
        weight_mem[16'h364B] <= 254;
        weight_mem[16'h364C] <= 17;
        weight_mem[16'h364D] <= 16;
        weight_mem[16'h364E] <= 22;
        weight_mem[16'h364F] <= 19;
        weight_mem[16'h3650] <= 23;
        weight_mem[16'h3651] <= 3;
        weight_mem[16'h3652] <= 5;
        weight_mem[16'h3653] <= 0;
        weight_mem[16'h3654] <= 224;
        weight_mem[16'h3655] <= 225;
        weight_mem[16'h3656] <= 213;
        weight_mem[16'h3657] <= 225;
        weight_mem[16'h3658] <= 233;
        weight_mem[16'h3659] <= 253;
        weight_mem[16'h365A] <= 8;
        weight_mem[16'h365B] <= 252;
        weight_mem[16'h365C] <= 255;
        weight_mem[16'h365D] <= 9;
        weight_mem[16'h365E] <= 254;
        weight_mem[16'h365F] <= 0;
        weight_mem[16'h3660] <= 251;
        weight_mem[16'h3661] <= 249;
        weight_mem[16'h3662] <= 3;
        weight_mem[16'h3663] <= 16;
        weight_mem[16'h3664] <= 16;
        weight_mem[16'h3665] <= 28;
        weight_mem[16'h3666] <= 20;
        weight_mem[16'h3667] <= 31;
        weight_mem[16'h3668] <= 48;
        weight_mem[16'h3669] <= 40;
        weight_mem[16'h366A] <= 36;
        weight_mem[16'h366B] <= 36;
        weight_mem[16'h366C] <= 7;
        weight_mem[16'h366D] <= 7;
        weight_mem[16'h366E] <= 8;
        weight_mem[16'h366F] <= 0;
        weight_mem[16'h3670] <= 15;
        weight_mem[16'h3671] <= 24;
        weight_mem[16'h3672] <= 15;
        weight_mem[16'h3673] <= 255;
        weight_mem[16'h3674] <= 1;
        weight_mem[16'h3675] <= 2;
        weight_mem[16'h3676] <= 251;
        weight_mem[16'h3677] <= 2;
        weight_mem[16'h3678] <= 4;
        weight_mem[16'h3679] <= 5;
        weight_mem[16'h367A] <= 11;
        weight_mem[16'h367B] <= 9;
        weight_mem[16'h367C] <= 33;
        weight_mem[16'h367D] <= 49;
        weight_mem[16'h367E] <= 40;
        weight_mem[16'h367F] <= 41;
        weight_mem[16'h3680] <= 32;
        weight_mem[16'h3681] <= 20;
        weight_mem[16'h3682] <= 30;
        weight_mem[16'h3683] <= 12;
        weight_mem[16'h3684] <= 14;
        weight_mem[16'h3685] <= 11;
        weight_mem[16'h3686] <= 244;
        weight_mem[16'h3687] <= 255;
        weight_mem[16'h3688] <= 18;
        weight_mem[16'h3689] <= 13;
        weight_mem[16'h368A] <= 12;
        weight_mem[16'h368B] <= 2;
        weight_mem[16'h368C] <= 253;
        weight_mem[16'h368D] <= 6;
        weight_mem[16'h368E] <= 8;
        weight_mem[16'h368F] <= 252;
        weight_mem[16'h3690] <= 4;
        weight_mem[16'h3691] <= 249;
        weight_mem[16'h3692] <= 11;
        weight_mem[16'h3693] <= 14;
        weight_mem[16'h3694] <= 32;
        weight_mem[16'h3695] <= 35;
        weight_mem[16'h3696] <= 38;
        weight_mem[16'h3697] <= 25;
        weight_mem[16'h3698] <= 14;
        weight_mem[16'h3699] <= 10;
        weight_mem[16'h369A] <= 10;
        weight_mem[16'h369B] <= 28;
        weight_mem[16'h369C] <= 58;
        weight_mem[16'h369D] <= 58;
        weight_mem[16'h369E] <= 8;
        weight_mem[16'h369F] <= 252;
        weight_mem[16'h36A0] <= 245;
        weight_mem[16'h36A1] <= 245;
        weight_mem[16'h36A2] <= 11;
        weight_mem[16'h36A3] <= 1;
        weight_mem[16'h36A4] <= 9;
        weight_mem[16'h36A5] <= 7;
        weight_mem[16'h36A6] <= 2;
        weight_mem[16'h36A7] <= 250;
        weight_mem[16'h36A8] <= 254;
        weight_mem[16'h36A9] <= 13;
        weight_mem[16'h36AA] <= 6;
        weight_mem[16'h36AB] <= 27;
        weight_mem[16'h36AC] <= 16;
        weight_mem[16'h36AD] <= 5;
        weight_mem[16'h36AE] <= 3;
        weight_mem[16'h36AF] <= 245;
        weight_mem[16'h36B0] <= 250;
        weight_mem[16'h36B1] <= 11;
        weight_mem[16'h36B2] <= 11;
        weight_mem[16'h36B3] <= 51;
        weight_mem[16'h36B4] <= 127;
        weight_mem[16'h36B5] <= 109;
        weight_mem[16'h36B6] <= 56;
        weight_mem[16'h36B7] <= 40;
        weight_mem[16'h36B8] <= 3;
        weight_mem[16'h36B9] <= 252;
        weight_mem[16'h36BA] <= 232;
        weight_mem[16'h36BB] <= 239;
        weight_mem[16'h36BC] <= 245;
        weight_mem[16'h36BD] <= 1;
        weight_mem[16'h36BE] <= 11;
        weight_mem[16'h36BF] <= 12;
        weight_mem[16'h36C0] <= 8;
        weight_mem[16'h36C1] <= 250;
        weight_mem[16'h36C2] <= 8;
        weight_mem[16'h36C3] <= 8;
        weight_mem[16'h36C4] <= 250;
        weight_mem[16'h36C5] <= 227;
        weight_mem[16'h36C6] <= 220;
        weight_mem[16'h36C7] <= 215;
        weight_mem[16'h36C8] <= 226;
        weight_mem[16'h36C9] <= 199;
        weight_mem[16'h36CA] <= 209;
        weight_mem[16'h36CB] <= 12;
        weight_mem[16'h36CC] <= 87;
        weight_mem[16'h36CD] <= 59;
        weight_mem[16'h36CE] <= 37;
        weight_mem[16'h36CF] <= 6;
        weight_mem[16'h36D0] <= 241;
        weight_mem[16'h36D1] <= 242;
        weight_mem[16'h36D2] <= 220;
        weight_mem[16'h36D3] <= 211;
        weight_mem[16'h36D4] <= 217;
        weight_mem[16'h36D5] <= 253;
        weight_mem[16'h36D6] <= 16;
        weight_mem[16'h36D7] <= 252;
        weight_mem[16'h36D8] <= 11;
        weight_mem[16'h36D9] <= 9;
        weight_mem[16'h36DA] <= 11;
        weight_mem[16'h36DB] <= 248;
        weight_mem[16'h36DC] <= 238;
        weight_mem[16'h36DD] <= 201;
        weight_mem[16'h36DE] <= 169;
        weight_mem[16'h36DF] <= 190;
        weight_mem[16'h36E0] <= 172;
        weight_mem[16'h36E1] <= 154;
        weight_mem[16'h36E2] <= 161;
        weight_mem[16'h36E3] <= 1;
        weight_mem[16'h36E4] <= 34;
        weight_mem[16'h36E5] <= 16;
        weight_mem[16'h36E6] <= 247;
        weight_mem[16'h36E7] <= 242;
        weight_mem[16'h36E8] <= 240;
        weight_mem[16'h36E9] <= 0;
        weight_mem[16'h36EA] <= 230;
        weight_mem[16'h36EB] <= 213;
        weight_mem[16'h36EC] <= 205;
        weight_mem[16'h36ED] <= 254;
        weight_mem[16'h36EE] <= 8;
        weight_mem[16'h36EF] <= 9;
        weight_mem[16'h36F0] <= 13;
        weight_mem[16'h36F1] <= 251;
        weight_mem[16'h36F2] <= 9;
        weight_mem[16'h36F3] <= 243;
        weight_mem[16'h36F4] <= 222;
        weight_mem[16'h36F5] <= 186;
        weight_mem[16'h36F6] <= 176;
        weight_mem[16'h36F7] <= 178;
        weight_mem[16'h36F8] <= 175;
        weight_mem[16'h36F9] <= 172;
        weight_mem[16'h36FA] <= 202;
        weight_mem[16'h36FB] <= 255;
        weight_mem[16'h36FC] <= 4;
        weight_mem[16'h36FD] <= 228;
        weight_mem[16'h36FE] <= 212;
        weight_mem[16'h36FF] <= 204;
        weight_mem[16'h3700] <= 231;
        weight_mem[16'h3701] <= 249;
        weight_mem[16'h3702] <= 228;
        weight_mem[16'h3703] <= 221;
        weight_mem[16'h3704] <= 233;
        weight_mem[16'h3705] <= 255;
        weight_mem[16'h3706] <= 0;
        weight_mem[16'h3707] <= 11;
        weight_mem[16'h3708] <= 9;
        weight_mem[16'h3709] <= 8;
        weight_mem[16'h370A] <= 253;
        weight_mem[16'h370B] <= 11;
        weight_mem[16'h370C] <= 225;
        weight_mem[16'h370D] <= 197;
        weight_mem[16'h370E] <= 188;
        weight_mem[16'h370F] <= 192;
        weight_mem[16'h3710] <= 187;
        weight_mem[16'h3711] <= 195;
        weight_mem[16'h3712] <= 228;
        weight_mem[16'h3713] <= 6;
        weight_mem[16'h3714] <= 11;
        weight_mem[16'h3715] <= 243;
        weight_mem[16'h3716] <= 203;
        weight_mem[16'h3717] <= 223;
        weight_mem[16'h3718] <= 225;
        weight_mem[16'h3719] <= 225;
        weight_mem[16'h371A] <= 219;
        weight_mem[16'h371B] <= 235;
        weight_mem[16'h371C] <= 252;
        weight_mem[16'h371D] <= 249;
        weight_mem[16'h371E] <= 12;
        weight_mem[16'h371F] <= 7;
        weight_mem[16'h3720] <= 247;
        weight_mem[16'h3721] <= 253;
        weight_mem[16'h3722] <= 13;
        weight_mem[16'h3723] <= 9;
        weight_mem[16'h3724] <= 0;
        weight_mem[16'h3725] <= 227;
        weight_mem[16'h3726] <= 218;
        weight_mem[16'h3727] <= 236;
        weight_mem[16'h3728] <= 225;
        weight_mem[16'h3729] <= 238;
        weight_mem[16'h372A] <= 250;
        weight_mem[16'h372B] <= 22;
        weight_mem[16'h372C] <= 15;
        weight_mem[16'h372D] <= 253;
        weight_mem[16'h372E] <= 249;
        weight_mem[16'h372F] <= 251;
        weight_mem[16'h3730] <= 247;
        weight_mem[16'h3731] <= 242;
        weight_mem[16'h3732] <= 242;
        weight_mem[16'h3733] <= 249;
        weight_mem[16'h3734] <= 10;
        weight_mem[16'h3735] <= 10;
        weight_mem[16'h3736] <= 14;
        weight_mem[16'h3737] <= 7;
        weight_mem[16'h3738] <= 4;
        weight_mem[16'h3739] <= 11;
        weight_mem[16'h373A] <= 12;
        weight_mem[16'h373B] <= 250;
        weight_mem[16'h373C] <= 246;
        weight_mem[16'h373D] <= 254;
        weight_mem[16'h373E] <= 251;
        weight_mem[16'h373F] <= 1;
        weight_mem[16'h3740] <= 0;
        weight_mem[16'h3741] <= 247;
        weight_mem[16'h3742] <= 224;
        weight_mem[16'h3743] <= 250;
        weight_mem[16'h3744] <= 2;
        weight_mem[16'h3745] <= 0;
        weight_mem[16'h3746] <= 12;
        weight_mem[16'h3747] <= 5;
        weight_mem[16'h3748] <= 250;
        weight_mem[16'h3749] <= 0;
        weight_mem[16'h374A] <= 243;
        weight_mem[16'h374B] <= 255;
        weight_mem[16'h374C] <= 6;
        weight_mem[16'h374D] <= 251;
        weight_mem[16'h374E] <= 249;
        weight_mem[16'h374F] <= 13;
        weight_mem[16'h3750] <= 8;
        weight_mem[16'h3751] <= 11;
        weight_mem[16'h3752] <= 7;
        weight_mem[16'h3753] <= 10;
        weight_mem[16'h3754] <= 18;
        weight_mem[16'h3755] <= 17;
        weight_mem[16'h3756] <= 4;
        weight_mem[16'h3757] <= 2;
        weight_mem[16'h3758] <= 235;
        weight_mem[16'h3759] <= 229;
        weight_mem[16'h375A] <= 219;
        weight_mem[16'h375B] <= 221;
        weight_mem[16'h375C] <= 243;
        weight_mem[16'h375D] <= 243;
        weight_mem[16'h375E] <= 6;
        weight_mem[16'h375F] <= 13;
        weight_mem[16'h3760] <= 7;
        weight_mem[16'h3761] <= 9;
        weight_mem[16'h3762] <= 252;
        weight_mem[16'h3763] <= 253;
        weight_mem[16'h3764] <= 15;
        weight_mem[16'h3765] <= 3;
        weight_mem[16'h3766] <= 11;
        weight_mem[16'h3767] <= 11;
        weight_mem[16'h3768] <= 3;
        weight_mem[16'h3769] <= 253;
        weight_mem[16'h376A] <= 6;
        weight_mem[16'h376B] <= 11;
        weight_mem[16'h376C] <= 8;
        weight_mem[16'h376D] <= 30;
        weight_mem[16'h376E] <= 17;
        weight_mem[16'h376F] <= 17;
        weight_mem[16'h3770] <= 24;
        weight_mem[16'h3771] <= 16;
        weight_mem[16'h3772] <= 9;
        weight_mem[16'h3773] <= 10;
        weight_mem[16'h3774] <= 13;
        weight_mem[16'h3775] <= 28;
        weight_mem[16'h3776] <= 38;
        weight_mem[16'h3777] <= 18;
        weight_mem[16'h3778] <= 8;
        weight_mem[16'h3779] <= 8;
        weight_mem[16'h377A] <= 6;
        weight_mem[16'h377B] <= 248;
        weight_mem[16'h377C] <= 11;
        weight_mem[16'h377D] <= 248;
        weight_mem[16'h377E] <= 7;
        weight_mem[16'h377F] <= 7;
        weight_mem[16'h3780] <= 250;
        weight_mem[16'h3781] <= 9;
        weight_mem[16'h3782] <= 252;
        weight_mem[16'h3783] <= 6;
        weight_mem[16'h3784] <= 2;
        weight_mem[16'h3785] <= 8;
        weight_mem[16'h3786] <= 13;
        weight_mem[16'h3787] <= 35;
        weight_mem[16'h3788] <= 45;
        weight_mem[16'h3789] <= 36;
        weight_mem[16'h378A] <= 46;
        weight_mem[16'h378B] <= 36;
        weight_mem[16'h378C] <= 38;
        weight_mem[16'h378D] <= 45;
        weight_mem[16'h378E] <= 40;
        weight_mem[16'h378F] <= 33;
        weight_mem[16'h3790] <= 28;
        weight_mem[16'h3791] <= 16;
        weight_mem[16'h3792] <= 7;
        weight_mem[16'h3793] <= 248;
        weight_mem[16'h3794] <= 5;
        weight_mem[16'h3795] <= 254;
        weight_mem[16'h3796] <= 5;
        weight_mem[16'h3797] <= 252;
        weight_mem[16'h3798] <= 2;
        weight_mem[16'h3799] <= 12;
        weight_mem[16'h379A] <= 252;
        weight_mem[16'h379B] <= 252;
        weight_mem[16'h379C] <= 254;
        weight_mem[16'h379D] <= 0;
        weight_mem[16'h379E] <= 251;
        weight_mem[16'h379F] <= 18;
        weight_mem[16'h37A0] <= 0;
        weight_mem[16'h37A1] <= 4;
        weight_mem[16'h37A2] <= 254;
        weight_mem[16'h37A3] <= 6;
        weight_mem[16'h37A4] <= 17;
        weight_mem[16'h37A5] <= 10;
        weight_mem[16'h37A6] <= 9;
        weight_mem[16'h37A7] <= 3;
        weight_mem[16'h37A8] <= 15;
        weight_mem[16'h37A9] <= 253;
        weight_mem[16'h37AA] <= 12;
        weight_mem[16'h37AB] <= 250;
        weight_mem[16'h37AC] <= 1;
        weight_mem[16'h37AD] <= 8;
        weight_mem[16'h37AE] <= 6;
        weight_mem[16'h37AF] <= 252;

        // layer 1 neuron 28
        weight_mem[16'h3800] <= 0;
        weight_mem[16'h3801] <= 0;
        weight_mem[16'h3802] <= 0;
        weight_mem[16'h3803] <= 0;
        weight_mem[16'h3804] <= 0;
        weight_mem[16'h3805] <= 0;
        weight_mem[16'h3806] <= 0;
        weight_mem[16'h3807] <= 0;
        weight_mem[16'h3808] <= 0;
        weight_mem[16'h3809] <= 0;
        weight_mem[16'h380A] <= 0;
        weight_mem[16'h380B] <= 0;
        weight_mem[16'h380C] <= 0;
        weight_mem[16'h380D] <= 0;
        weight_mem[16'h380E] <= 0;
        weight_mem[16'h380F] <= 0;
        weight_mem[16'h3810] <= 0;
        weight_mem[16'h3811] <= 0;
        weight_mem[16'h3812] <= 0;
        weight_mem[16'h3813] <= 0;
        weight_mem[16'h3814] <= 0;
        weight_mem[16'h3815] <= 0;
        weight_mem[16'h3816] <= 0;
        weight_mem[16'h3817] <= 0;
        weight_mem[16'h3818] <= 0;
        weight_mem[16'h3819] <= 0;
        weight_mem[16'h381A] <= 0;
        weight_mem[16'h381B] <= 0;
        weight_mem[16'h381C] <= 0;
        weight_mem[16'h381D] <= 0;
        weight_mem[16'h381E] <= 0;
        weight_mem[16'h381F] <= 0;
        weight_mem[16'h3820] <= 0;
        weight_mem[16'h3821] <= 0;
        weight_mem[16'h3822] <= 0;
        weight_mem[16'h3823] <= 0;
        weight_mem[16'h3824] <= 0;
        weight_mem[16'h3825] <= 0;
        weight_mem[16'h3826] <= 0;
        weight_mem[16'h3827] <= 0;
        weight_mem[16'h3828] <= 0;
        weight_mem[16'h3829] <= 0;
        weight_mem[16'h382A] <= 0;
        weight_mem[16'h382B] <= 0;
        weight_mem[16'h382C] <= 0;
        weight_mem[16'h382D] <= 0;
        weight_mem[16'h382E] <= 0;
        weight_mem[16'h382F] <= 0;
        weight_mem[16'h3830] <= 0;
        weight_mem[16'h3831] <= 0;
        weight_mem[16'h3832] <= 0;
        weight_mem[16'h3833] <= 0;
        weight_mem[16'h3834] <= 0;
        weight_mem[16'h3835] <= 0;
        weight_mem[16'h3836] <= 0;
        weight_mem[16'h3837] <= 0;
        weight_mem[16'h3838] <= 0;
        weight_mem[16'h3839] <= 0;
        weight_mem[16'h383A] <= 0;
        weight_mem[16'h383B] <= 0;
        weight_mem[16'h383C] <= 0;
        weight_mem[16'h383D] <= 0;
        weight_mem[16'h383E] <= 0;
        weight_mem[16'h383F] <= 0;
        weight_mem[16'h3840] <= 0;
        weight_mem[16'h3841] <= 0;
        weight_mem[16'h3842] <= 0;
        weight_mem[16'h3843] <= 0;
        weight_mem[16'h3844] <= 0;
        weight_mem[16'h3845] <= 0;
        weight_mem[16'h3846] <= 0;
        weight_mem[16'h3847] <= 0;
        weight_mem[16'h3848] <= 0;
        weight_mem[16'h3849] <= 0;
        weight_mem[16'h384A] <= 0;
        weight_mem[16'h384B] <= 0;
        weight_mem[16'h384C] <= 0;
        weight_mem[16'h384D] <= 0;
        weight_mem[16'h384E] <= 0;
        weight_mem[16'h384F] <= 0;
        weight_mem[16'h3850] <= 0;
        weight_mem[16'h3851] <= 0;
        weight_mem[16'h3852] <= 0;
        weight_mem[16'h3853] <= 0;
        weight_mem[16'h3854] <= 0;
        weight_mem[16'h3855] <= 0;
        weight_mem[16'h3856] <= 0;
        weight_mem[16'h3857] <= 0;
        weight_mem[16'h3858] <= 0;
        weight_mem[16'h3859] <= 0;
        weight_mem[16'h385A] <= 0;
        weight_mem[16'h385B] <= 0;
        weight_mem[16'h385C] <= 0;
        weight_mem[16'h385D] <= 0;
        weight_mem[16'h385E] <= 0;
        weight_mem[16'h385F] <= 0;
        weight_mem[16'h3860] <= 0;
        weight_mem[16'h3861] <= 0;
        weight_mem[16'h3862] <= 0;
        weight_mem[16'h3863] <= 0;
        weight_mem[16'h3864] <= 0;
        weight_mem[16'h3865] <= 0;
        weight_mem[16'h3866] <= 0;
        weight_mem[16'h3867] <= 0;
        weight_mem[16'h3868] <= 0;
        weight_mem[16'h3869] <= 0;
        weight_mem[16'h386A] <= 0;
        weight_mem[16'h386B] <= 0;
        weight_mem[16'h386C] <= 0;
        weight_mem[16'h386D] <= 0;
        weight_mem[16'h386E] <= 0;
        weight_mem[16'h386F] <= 0;
        weight_mem[16'h3870] <= 0;
        weight_mem[16'h3871] <= 0;
        weight_mem[16'h3872] <= 0;
        weight_mem[16'h3873] <= 0;
        weight_mem[16'h3874] <= 0;
        weight_mem[16'h3875] <= 0;
        weight_mem[16'h3876] <= 0;
        weight_mem[16'h3877] <= 0;
        weight_mem[16'h3878] <= 0;
        weight_mem[16'h3879] <= 0;
        weight_mem[16'h387A] <= 0;
        weight_mem[16'h387B] <= 0;
        weight_mem[16'h387C] <= 0;
        weight_mem[16'h387D] <= 0;
        weight_mem[16'h387E] <= 0;
        weight_mem[16'h387F] <= 0;
        weight_mem[16'h3880] <= 0;
        weight_mem[16'h3881] <= 0;
        weight_mem[16'h3882] <= 0;
        weight_mem[16'h3883] <= 0;
        weight_mem[16'h3884] <= 0;
        weight_mem[16'h3885] <= 0;
        weight_mem[16'h3886] <= 0;
        weight_mem[16'h3887] <= 0;
        weight_mem[16'h3888] <= 0;
        weight_mem[16'h3889] <= 0;
        weight_mem[16'h388A] <= 0;
        weight_mem[16'h388B] <= 0;
        weight_mem[16'h388C] <= 0;
        weight_mem[16'h388D] <= 0;
        weight_mem[16'h388E] <= 0;
        weight_mem[16'h388F] <= 0;
        weight_mem[16'h3890] <= 0;
        weight_mem[16'h3891] <= 0;
        weight_mem[16'h3892] <= 0;
        weight_mem[16'h3893] <= 0;
        weight_mem[16'h3894] <= 0;
        weight_mem[16'h3895] <= 0;
        weight_mem[16'h3896] <= 0;
        weight_mem[16'h3897] <= 0;
        weight_mem[16'h3898] <= 0;
        weight_mem[16'h3899] <= 0;
        weight_mem[16'h389A] <= 0;
        weight_mem[16'h389B] <= 0;
        weight_mem[16'h389C] <= 0;
        weight_mem[16'h389D] <= 0;
        weight_mem[16'h389E] <= 0;
        weight_mem[16'h389F] <= 0;
        weight_mem[16'h38A0] <= 0;
        weight_mem[16'h38A1] <= 0;
        weight_mem[16'h38A2] <= 0;
        weight_mem[16'h38A3] <= 0;
        weight_mem[16'h38A4] <= 0;
        weight_mem[16'h38A5] <= 0;
        weight_mem[16'h38A6] <= 0;
        weight_mem[16'h38A7] <= 0;
        weight_mem[16'h38A8] <= 0;
        weight_mem[16'h38A9] <= 0;
        weight_mem[16'h38AA] <= 0;
        weight_mem[16'h38AB] <= 0;
        weight_mem[16'h38AC] <= 0;
        weight_mem[16'h38AD] <= 0;
        weight_mem[16'h38AE] <= 0;
        weight_mem[16'h38AF] <= 0;
        weight_mem[16'h38B0] <= 0;
        weight_mem[16'h38B1] <= 0;
        weight_mem[16'h38B2] <= 0;
        weight_mem[16'h38B3] <= 0;
        weight_mem[16'h38B4] <= 0;
        weight_mem[16'h38B5] <= 0;
        weight_mem[16'h38B6] <= 0;
        weight_mem[16'h38B7] <= 0;
        weight_mem[16'h38B8] <= 0;
        weight_mem[16'h38B9] <= 0;
        weight_mem[16'h38BA] <= 0;
        weight_mem[16'h38BB] <= 0;
        weight_mem[16'h38BC] <= 0;
        weight_mem[16'h38BD] <= 0;
        weight_mem[16'h38BE] <= 0;
        weight_mem[16'h38BF] <= 0;
        weight_mem[16'h38C0] <= 0;
        weight_mem[16'h38C1] <= 0;
        weight_mem[16'h38C2] <= 0;
        weight_mem[16'h38C3] <= 0;
        weight_mem[16'h38C4] <= 0;
        weight_mem[16'h38C5] <= 0;
        weight_mem[16'h38C6] <= 0;
        weight_mem[16'h38C7] <= 0;
        weight_mem[16'h38C8] <= 0;
        weight_mem[16'h38C9] <= 0;
        weight_mem[16'h38CA] <= 0;
        weight_mem[16'h38CB] <= 0;
        weight_mem[16'h38CC] <= 0;
        weight_mem[16'h38CD] <= 0;
        weight_mem[16'h38CE] <= 0;
        weight_mem[16'h38CF] <= 0;
        weight_mem[16'h38D0] <= 0;
        weight_mem[16'h38D1] <= 0;
        weight_mem[16'h38D2] <= 0;
        weight_mem[16'h38D3] <= 0;
        weight_mem[16'h38D4] <= 0;
        weight_mem[16'h38D5] <= 0;
        weight_mem[16'h38D6] <= 0;
        weight_mem[16'h38D7] <= 0;
        weight_mem[16'h38D8] <= 0;
        weight_mem[16'h38D9] <= 0;
        weight_mem[16'h38DA] <= 0;
        weight_mem[16'h38DB] <= 0;
        weight_mem[16'h38DC] <= 0;
        weight_mem[16'h38DD] <= 0;
        weight_mem[16'h38DE] <= 0;
        weight_mem[16'h38DF] <= 0;
        weight_mem[16'h38E0] <= 0;
        weight_mem[16'h38E1] <= 0;
        weight_mem[16'h38E2] <= 0;
        weight_mem[16'h38E3] <= 0;
        weight_mem[16'h38E4] <= 0;
        weight_mem[16'h38E5] <= 0;
        weight_mem[16'h38E6] <= 0;
        weight_mem[16'h38E7] <= 0;
        weight_mem[16'h38E8] <= 0;
        weight_mem[16'h38E9] <= 0;
        weight_mem[16'h38EA] <= 0;
        weight_mem[16'h38EB] <= 0;
        weight_mem[16'h38EC] <= 0;
        weight_mem[16'h38ED] <= 0;
        weight_mem[16'h38EE] <= 0;
        weight_mem[16'h38EF] <= 0;
        weight_mem[16'h38F0] <= 0;
        weight_mem[16'h38F1] <= 0;
        weight_mem[16'h38F2] <= 0;
        weight_mem[16'h38F3] <= 0;
        weight_mem[16'h38F4] <= 0;
        weight_mem[16'h38F5] <= 0;
        weight_mem[16'h38F6] <= 0;
        weight_mem[16'h38F7] <= 0;
        weight_mem[16'h38F8] <= 0;
        weight_mem[16'h38F9] <= 0;
        weight_mem[16'h38FA] <= 0;
        weight_mem[16'h38FB] <= 0;
        weight_mem[16'h38FC] <= 0;
        weight_mem[16'h38FD] <= 0;
        weight_mem[16'h38FE] <= 0;
        weight_mem[16'h38FF] <= 0;
        weight_mem[16'h3900] <= 0;
        weight_mem[16'h3901] <= 0;
        weight_mem[16'h3902] <= 0;
        weight_mem[16'h3903] <= 0;
        weight_mem[16'h3904] <= 0;
        weight_mem[16'h3905] <= 0;
        weight_mem[16'h3906] <= 0;
        weight_mem[16'h3907] <= 0;
        weight_mem[16'h3908] <= 0;
        weight_mem[16'h3909] <= 0;
        weight_mem[16'h390A] <= 0;
        weight_mem[16'h390B] <= 0;
        weight_mem[16'h390C] <= 0;
        weight_mem[16'h390D] <= 0;
        weight_mem[16'h390E] <= 0;
        weight_mem[16'h390F] <= 0;
        weight_mem[16'h3910] <= 0;
        weight_mem[16'h3911] <= 0;
        weight_mem[16'h3912] <= 0;
        weight_mem[16'h3913] <= 0;
        weight_mem[16'h3914] <= 0;
        weight_mem[16'h3915] <= 0;
        weight_mem[16'h3916] <= 0;
        weight_mem[16'h3917] <= 0;
        weight_mem[16'h3918] <= 0;
        weight_mem[16'h3919] <= 0;
        weight_mem[16'h391A] <= 0;
        weight_mem[16'h391B] <= 0;
        weight_mem[16'h391C] <= 0;
        weight_mem[16'h391D] <= 0;
        weight_mem[16'h391E] <= 0;
        weight_mem[16'h391F] <= 0;
        weight_mem[16'h3920] <= 0;
        weight_mem[16'h3921] <= 0;
        weight_mem[16'h3922] <= 0;
        weight_mem[16'h3923] <= 0;
        weight_mem[16'h3924] <= 0;
        weight_mem[16'h3925] <= 0;
        weight_mem[16'h3926] <= 0;
        weight_mem[16'h3927] <= 0;
        weight_mem[16'h3928] <= 0;
        weight_mem[16'h3929] <= 0;
        weight_mem[16'h392A] <= 0;
        weight_mem[16'h392B] <= 0;
        weight_mem[16'h392C] <= 0;
        weight_mem[16'h392D] <= 0;
        weight_mem[16'h392E] <= 0;
        weight_mem[16'h392F] <= 0;
        weight_mem[16'h3930] <= 0;
        weight_mem[16'h3931] <= 0;
        weight_mem[16'h3932] <= 0;
        weight_mem[16'h3933] <= 0;
        weight_mem[16'h3934] <= 0;
        weight_mem[16'h3935] <= 0;
        weight_mem[16'h3936] <= 0;
        weight_mem[16'h3937] <= 0;
        weight_mem[16'h3938] <= 0;
        weight_mem[16'h3939] <= 0;
        weight_mem[16'h393A] <= 0;
        weight_mem[16'h393B] <= 0;
        weight_mem[16'h393C] <= 0;
        weight_mem[16'h393D] <= 0;
        weight_mem[16'h393E] <= 0;
        weight_mem[16'h393F] <= 0;
        weight_mem[16'h3940] <= 0;
        weight_mem[16'h3941] <= 0;
        weight_mem[16'h3942] <= 0;
        weight_mem[16'h3943] <= 0;
        weight_mem[16'h3944] <= 0;
        weight_mem[16'h3945] <= 0;
        weight_mem[16'h3946] <= 0;
        weight_mem[16'h3947] <= 0;
        weight_mem[16'h3948] <= 0;
        weight_mem[16'h3949] <= 0;
        weight_mem[16'h394A] <= 0;
        weight_mem[16'h394B] <= 0;
        weight_mem[16'h394C] <= 0;
        weight_mem[16'h394D] <= 0;
        weight_mem[16'h394E] <= 0;
        weight_mem[16'h394F] <= 0;
        weight_mem[16'h3950] <= 0;
        weight_mem[16'h3951] <= 0;
        weight_mem[16'h3952] <= 0;
        weight_mem[16'h3953] <= 0;
        weight_mem[16'h3954] <= 0;
        weight_mem[16'h3955] <= 0;
        weight_mem[16'h3956] <= 0;
        weight_mem[16'h3957] <= 0;
        weight_mem[16'h3958] <= 0;
        weight_mem[16'h3959] <= 0;
        weight_mem[16'h395A] <= 0;
        weight_mem[16'h395B] <= 0;
        weight_mem[16'h395C] <= 0;
        weight_mem[16'h395D] <= 0;
        weight_mem[16'h395E] <= 0;
        weight_mem[16'h395F] <= 0;
        weight_mem[16'h3960] <= 0;
        weight_mem[16'h3961] <= 0;
        weight_mem[16'h3962] <= 0;
        weight_mem[16'h3963] <= 0;
        weight_mem[16'h3964] <= 0;
        weight_mem[16'h3965] <= 0;
        weight_mem[16'h3966] <= 0;
        weight_mem[16'h3967] <= 0;
        weight_mem[16'h3968] <= 0;
        weight_mem[16'h3969] <= 0;
        weight_mem[16'h396A] <= 0;
        weight_mem[16'h396B] <= 0;
        weight_mem[16'h396C] <= 0;
        weight_mem[16'h396D] <= 0;
        weight_mem[16'h396E] <= 0;
        weight_mem[16'h396F] <= 0;
        weight_mem[16'h3970] <= 0;
        weight_mem[16'h3971] <= 0;
        weight_mem[16'h3972] <= 0;
        weight_mem[16'h3973] <= 0;
        weight_mem[16'h3974] <= 0;
        weight_mem[16'h3975] <= 0;
        weight_mem[16'h3976] <= 0;
        weight_mem[16'h3977] <= 0;
        weight_mem[16'h3978] <= 0;
        weight_mem[16'h3979] <= 0;
        weight_mem[16'h397A] <= 0;
        weight_mem[16'h397B] <= 0;
        weight_mem[16'h397C] <= 0;
        weight_mem[16'h397D] <= 0;
        weight_mem[16'h397E] <= 0;
        weight_mem[16'h397F] <= 0;
        weight_mem[16'h3980] <= 0;
        weight_mem[16'h3981] <= 0;
        weight_mem[16'h3982] <= 0;
        weight_mem[16'h3983] <= 0;
        weight_mem[16'h3984] <= 0;
        weight_mem[16'h3985] <= 0;
        weight_mem[16'h3986] <= 0;
        weight_mem[16'h3987] <= 0;
        weight_mem[16'h3988] <= 0;
        weight_mem[16'h3989] <= 0;
        weight_mem[16'h398A] <= 0;
        weight_mem[16'h398B] <= 0;
        weight_mem[16'h398C] <= 0;
        weight_mem[16'h398D] <= 0;
        weight_mem[16'h398E] <= 0;
        weight_mem[16'h398F] <= 0;
        weight_mem[16'h3990] <= 0;
        weight_mem[16'h3991] <= 0;
        weight_mem[16'h3992] <= 0;
        weight_mem[16'h3993] <= 0;
        weight_mem[16'h3994] <= 0;
        weight_mem[16'h3995] <= 0;
        weight_mem[16'h3996] <= 0;
        weight_mem[16'h3997] <= 0;
        weight_mem[16'h3998] <= 0;
        weight_mem[16'h3999] <= 0;
        weight_mem[16'h399A] <= 0;
        weight_mem[16'h399B] <= 0;
        weight_mem[16'h399C] <= 0;
        weight_mem[16'h399D] <= 0;
        weight_mem[16'h399E] <= 0;
        weight_mem[16'h399F] <= 0;
        weight_mem[16'h39A0] <= 0;
        weight_mem[16'h39A1] <= 0;
        weight_mem[16'h39A2] <= 0;
        weight_mem[16'h39A3] <= 0;
        weight_mem[16'h39A4] <= 0;
        weight_mem[16'h39A5] <= 0;
        weight_mem[16'h39A6] <= 0;
        weight_mem[16'h39A7] <= 0;
        weight_mem[16'h39A8] <= 0;
        weight_mem[16'h39A9] <= 0;
        weight_mem[16'h39AA] <= 0;
        weight_mem[16'h39AB] <= 0;
        weight_mem[16'h39AC] <= 0;
        weight_mem[16'h39AD] <= 0;
        weight_mem[16'h39AE] <= 0;
        weight_mem[16'h39AF] <= 0;

        // layer 1 neuron 29
        weight_mem[16'h3A00] <= 232;
        weight_mem[16'h3A01] <= 237;
        weight_mem[16'h3A02] <= 234;
        weight_mem[16'h3A03] <= 246;
        weight_mem[16'h3A04] <= 244;
        weight_mem[16'h3A05] <= 236;
        weight_mem[16'h3A06] <= 239;
        weight_mem[16'h3A07] <= 248;
        weight_mem[16'h3A08] <= 249;
        weight_mem[16'h3A09] <= 252;
        weight_mem[16'h3A0A] <= 245;
        weight_mem[16'h3A0B] <= 230;
        weight_mem[16'h3A0C] <= 234;
        weight_mem[16'h3A0D] <= 232;
        weight_mem[16'h3A0E] <= 245;
        weight_mem[16'h3A0F] <= 239;
        weight_mem[16'h3A10] <= 235;
        weight_mem[16'h3A11] <= 231;
        weight_mem[16'h3A12] <= 246;
        weight_mem[16'h3A13] <= 239;
        weight_mem[16'h3A14] <= 246;
        weight_mem[16'h3A15] <= 241;
        weight_mem[16'h3A16] <= 236;
        weight_mem[16'h3A17] <= 231;
        weight_mem[16'h3A18] <= 235;
        weight_mem[16'h3A19] <= 247;
        weight_mem[16'h3A1A] <= 235;
        weight_mem[16'h3A1B] <= 246;
        weight_mem[16'h3A1C] <= 243;
        weight_mem[16'h3A1D] <= 247;
        weight_mem[16'h3A1E] <= 239;
        weight_mem[16'h3A1F] <= 238;
        weight_mem[16'h3A20] <= 235;
        weight_mem[16'h3A21] <= 234;
        weight_mem[16'h3A22] <= 239;
        weight_mem[16'h3A23] <= 252;
        weight_mem[16'h3A24] <= 245;
        weight_mem[16'h3A25] <= 252;
        weight_mem[16'h3A26] <= 248;
        weight_mem[16'h3A27] <= 243;
        weight_mem[16'h3A28] <= 250;
        weight_mem[16'h3A29] <= 243;
        weight_mem[16'h3A2A] <= 246;
        weight_mem[16'h3A2B] <= 251;
        weight_mem[16'h3A2C] <= 250;
        weight_mem[16'h3A2D] <= 244;
        weight_mem[16'h3A2E] <= 242;
        weight_mem[16'h3A2F] <= 232;
        weight_mem[16'h3A30] <= 253;
        weight_mem[16'h3A31] <= 232;
        weight_mem[16'h3A32] <= 253;
        weight_mem[16'h3A33] <= 248;
        weight_mem[16'h3A34] <= 231;
        weight_mem[16'h3A35] <= 240;
        weight_mem[16'h3A36] <= 246;
        weight_mem[16'h3A37] <= 3;
        weight_mem[16'h3A38] <= 15;
        weight_mem[16'h3A39] <= 5;
        weight_mem[16'h3A3A] <= 15;
        weight_mem[16'h3A3B] <= 13;
        weight_mem[16'h3A3C] <= 3;
        weight_mem[16'h3A3D] <= 1;
        weight_mem[16'h3A3E] <= 248;
        weight_mem[16'h3A3F] <= 243;
        weight_mem[16'h3A40] <= 244;
        weight_mem[16'h3A41] <= 231;
        weight_mem[16'h3A42] <= 242;
        weight_mem[16'h3A43] <= 232;
        weight_mem[16'h3A44] <= 239;
        weight_mem[16'h3A45] <= 246;
        weight_mem[16'h3A46] <= 243;
        weight_mem[16'h3A47] <= 244;
        weight_mem[16'h3A48] <= 248;
        weight_mem[16'h3A49] <= 246;
        weight_mem[16'h3A4A] <= 242;
        weight_mem[16'h3A4B] <= 236;
        weight_mem[16'h3A4C] <= 255;
        weight_mem[16'h3A4D] <= 2;
        weight_mem[16'h3A4E] <= 22;
        weight_mem[16'h3A4F] <= 30;
        weight_mem[16'h3A50] <= 54;
        weight_mem[16'h3A51] <= 51;
        weight_mem[16'h3A52] <= 56;
        weight_mem[16'h3A53] <= 42;
        weight_mem[16'h3A54] <= 25;
        weight_mem[16'h3A55] <= 20;
        weight_mem[16'h3A56] <= 47;
        weight_mem[16'h3A57] <= 29;
        weight_mem[16'h3A58] <= 17;
        weight_mem[16'h3A59] <= 15;
        weight_mem[16'h3A5A] <= 234;
        weight_mem[16'h3A5B] <= 217;
        weight_mem[16'h3A5C] <= 225;
        weight_mem[16'h3A5D] <= 254;
        weight_mem[16'h3A5E] <= 234;
        weight_mem[16'h3A5F] <= 247;
        weight_mem[16'h3A60] <= 234;
        weight_mem[16'h3A61] <= 246;
        weight_mem[16'h3A62] <= 240;
        weight_mem[16'h3A63] <= 242;
        weight_mem[16'h3A64] <= 249;
        weight_mem[16'h3A65] <= 27;
        weight_mem[16'h3A66] <= 34;
        weight_mem[16'h3A67] <= 58;
        weight_mem[16'h3A68] <= 52;
        weight_mem[16'h3A69] <= 22;
        weight_mem[16'h3A6A] <= 11;
        weight_mem[16'h3A6B] <= 2;
        weight_mem[16'h3A6C] <= 240;
        weight_mem[16'h3A6D] <= 242;
        weight_mem[16'h3A6E] <= 251;
        weight_mem[16'h3A6F] <= 12;
        weight_mem[16'h3A70] <= 14;
        weight_mem[16'h3A71] <= 5;
        weight_mem[16'h3A72] <= 254;
        weight_mem[16'h3A73] <= 232;
        weight_mem[16'h3A74] <= 6;
        weight_mem[16'h3A75] <= 245;
        weight_mem[16'h3A76] <= 238;
        weight_mem[16'h3A77] <= 231;
        weight_mem[16'h3A78] <= 253;
        weight_mem[16'h3A79] <= 252;
        weight_mem[16'h3A7A] <= 250;
        weight_mem[16'h3A7B] <= 1;
        weight_mem[16'h3A7C] <= 17;
        weight_mem[16'h3A7D] <= 36;
        weight_mem[16'h3A7E] <= 38;
        weight_mem[16'h3A7F] <= 55;
        weight_mem[16'h3A80] <= 42;
        weight_mem[16'h3A81] <= 26;
        weight_mem[16'h3A82] <= 6;
        weight_mem[16'h3A83] <= 242;
        weight_mem[16'h3A84] <= 226;
        weight_mem[16'h3A85] <= 243;
        weight_mem[16'h3A86] <= 2;
        weight_mem[16'h3A87] <= 0;
        weight_mem[16'h3A88] <= 6;
        weight_mem[16'h3A89] <= 11;
        weight_mem[16'h3A8A] <= 20;
        weight_mem[16'h3A8B] <= 16;
        weight_mem[16'h3A8C] <= 28;
        weight_mem[16'h3A8D] <= 12;
        weight_mem[16'h3A8E] <= 250;
        weight_mem[16'h3A8F] <= 249;
        weight_mem[16'h3A90] <= 254;
        weight_mem[16'h3A91] <= 230;
        weight_mem[16'h3A92] <= 249;
        weight_mem[16'h3A93] <= 246;
        weight_mem[16'h3A94] <= 254;
        weight_mem[16'h3A95] <= 34;
        weight_mem[16'h3A96] <= 47;
        weight_mem[16'h3A97] <= 37;
        weight_mem[16'h3A98] <= 35;
        weight_mem[16'h3A99] <= 27;
        weight_mem[16'h3A9A] <= 7;
        weight_mem[16'h3A9B] <= 232;
        weight_mem[16'h3A9C] <= 200;
        weight_mem[16'h3A9D] <= 215;
        weight_mem[16'h3A9E] <= 19;
        weight_mem[16'h3A9F] <= 44;
        weight_mem[16'h3AA0] <= 40;
        weight_mem[16'h3AA1] <= 44;
        weight_mem[16'h3AA2] <= 24;
        weight_mem[16'h3AA3] <= 43;
        weight_mem[16'h3AA4] <= 45;
        weight_mem[16'h3AA5] <= 27;
        weight_mem[16'h3AA6] <= 0;
        weight_mem[16'h3AA7] <= 237;
        weight_mem[16'h3AA8] <= 237;
        weight_mem[16'h3AA9] <= 235;
        weight_mem[16'h3AAA] <= 238;
        weight_mem[16'h3AAB] <= 249;
        weight_mem[16'h3AAC] <= 5;
        weight_mem[16'h3AAD] <= 23;
        weight_mem[16'h3AAE] <= 15;
        weight_mem[16'h3AAF] <= 0;
        weight_mem[16'h3AB0] <= 242;
        weight_mem[16'h3AB1] <= 236;
        weight_mem[16'h3AB2] <= 225;
        weight_mem[16'h3AB3] <= 204;
        weight_mem[16'h3AB4] <= 167;
        weight_mem[16'h3AB5] <= 169;
        weight_mem[16'h3AB6] <= 8;
        weight_mem[16'h3AB7] <= 22;
        weight_mem[16'h3AB8] <= 11;
        weight_mem[16'h3AB9] <= 12;
        weight_mem[16'h3ABA] <= 15;
        weight_mem[16'h3ABB] <= 17;
        weight_mem[16'h3ABC] <= 12;
        weight_mem[16'h3ABD] <= 253;
        weight_mem[16'h3ABE] <= 249;
        weight_mem[16'h3ABF] <= 250;
        weight_mem[16'h3AC0] <= 238;
        weight_mem[16'h3AC1] <= 239;
        weight_mem[16'h3AC2] <= 244;
        weight_mem[16'h3AC3] <= 245;
        weight_mem[16'h3AC4] <= 236;
        weight_mem[16'h3AC5] <= 253;
        weight_mem[16'h3AC6] <= 243;
        weight_mem[16'h3AC7] <= 244;
        weight_mem[16'h3AC8] <= 212;
        weight_mem[16'h3AC9] <= 230;
        weight_mem[16'h3ACA] <= 224;
        weight_mem[16'h3ACB] <= 207;
        weight_mem[16'h3ACC] <= 129;
        weight_mem[16'h3ACD] <= 166;
        weight_mem[16'h3ACE] <= 229;
        weight_mem[16'h3ACF] <= 247;
        weight_mem[16'h3AD0] <= 1;
        weight_mem[16'h3AD1] <= 253;
        weight_mem[16'h3AD2] <= 12;
        weight_mem[16'h3AD3] <= 19;
        weight_mem[16'h3AD4] <= 22;
        weight_mem[16'h3AD5] <= 252;
        weight_mem[16'h3AD6] <= 254;
        weight_mem[16'h3AD7] <= 243;
        weight_mem[16'h3AD8] <= 234;
        weight_mem[16'h3AD9] <= 237;
        weight_mem[16'h3ADA] <= 241;
        weight_mem[16'h3ADB] <= 234;
        weight_mem[16'h3ADC] <= 248;
        weight_mem[16'h3ADD] <= 13;
        weight_mem[16'h3ADE] <= 10;
        weight_mem[16'h3ADF] <= 1;
        weight_mem[16'h3AE0] <= 244;
        weight_mem[16'h3AE1] <= 237;
        weight_mem[16'h3AE2] <= 238;
        weight_mem[16'h3AE3] <= 202;
        weight_mem[16'h3AE4] <= 167;
        weight_mem[16'h3AE5] <= 166;
        weight_mem[16'h3AE6] <= 223;
        weight_mem[16'h3AE7] <= 0;
        weight_mem[16'h3AE8] <= 13;
        weight_mem[16'h3AE9] <= 25;
        weight_mem[16'h3AEA] <= 6;
        weight_mem[16'h3AEB] <= 8;
        weight_mem[16'h3AEC] <= 14;
        weight_mem[16'h3AED] <= 254;
        weight_mem[16'h3AEE] <= 244;
        weight_mem[16'h3AEF] <= 240;
        weight_mem[16'h3AF0] <= 247;
        weight_mem[16'h3AF1] <= 238;
        weight_mem[16'h3AF2] <= 236;
        weight_mem[16'h3AF3] <= 252;
        weight_mem[16'h3AF4] <= 12;
        weight_mem[16'h3AF5] <= 44;
        weight_mem[16'h3AF6] <= 47;
        weight_mem[16'h3AF7] <= 24;
        weight_mem[16'h3AF8] <= 3;
        weight_mem[16'h3AF9] <= 240;
        weight_mem[16'h3AFA] <= 1;
        weight_mem[16'h3AFB] <= 233;
        weight_mem[16'h3AFC] <= 176;
        weight_mem[16'h3AFD] <= 203;
        weight_mem[16'h3AFE] <= 8;
        weight_mem[16'h3AFF] <= 52;
        weight_mem[16'h3B00] <= 43;
        weight_mem[16'h3B01] <= 46;
        weight_mem[16'h3B02] <= 25;
        weight_mem[16'h3B03] <= 30;
        weight_mem[16'h3B04] <= 10;
        weight_mem[16'h3B05] <= 11;
        weight_mem[16'h3B06] <= 5;
        weight_mem[16'h3B07] <= 242;
        weight_mem[16'h3B08] <= 234;
        weight_mem[16'h3B09] <= 233;
        weight_mem[16'h3B0A] <= 237;
        weight_mem[16'h3B0B] <= 250;
        weight_mem[16'h3B0C] <= 20;
        weight_mem[16'h3B0D] <= 81;
        weight_mem[16'h3B0E] <= 88;
        weight_mem[16'h3B0F] <= 69;
        weight_mem[16'h3B10] <= 43;
        weight_mem[16'h3B11] <= 27;
        weight_mem[16'h3B12] <= 6;
        weight_mem[16'h3B13] <= 208;
        weight_mem[16'h3B14] <= 187;
        weight_mem[16'h3B15] <= 15;
        weight_mem[16'h3B16] <= 83;
        weight_mem[16'h3B17] <= 77;
        weight_mem[16'h3B18] <= 74;
        weight_mem[16'h3B19] <= 57;
        weight_mem[16'h3B1A] <= 45;
        weight_mem[16'h3B1B] <= 55;
        weight_mem[16'h3B1C] <= 33;
        weight_mem[16'h3B1D] <= 22;
        weight_mem[16'h3B1E] <= 4;
        weight_mem[16'h3B1F] <= 249;
        weight_mem[16'h3B20] <= 245;
        weight_mem[16'h3B21] <= 253;
        weight_mem[16'h3B22] <= 252;
        weight_mem[16'h3B23] <= 251;
        weight_mem[16'h3B24] <= 42;
        weight_mem[16'h3B25] <= 65;
        weight_mem[16'h3B26] <= 99;
        weight_mem[16'h3B27] <= 92;
        weight_mem[16'h3B28] <= 53;
        weight_mem[16'h3B29] <= 22;
        weight_mem[16'h3B2A] <= 253;
        weight_mem[16'h3B2B] <= 216;
        weight_mem[16'h3B2C] <= 243;
        weight_mem[16'h3B2D] <= 44;
        weight_mem[16'h3B2E] <= 72;
        weight_mem[16'h3B2F] <= 65;
        weight_mem[16'h3B30] <= 69;
        weight_mem[16'h3B31] <= 54;
        weight_mem[16'h3B32] <= 46;
        weight_mem[16'h3B33] <= 38;
        weight_mem[16'h3B34] <= 22;
        weight_mem[16'h3B35] <= 4;
        weight_mem[16'h3B36] <= 248;
        weight_mem[16'h3B37] <= 236;
        weight_mem[16'h3B38] <= 243;
        weight_mem[16'h3B39] <= 233;
        weight_mem[16'h3B3A] <= 245;
        weight_mem[16'h3B3B] <= 10;
        weight_mem[16'h3B3C] <= 22;
        weight_mem[16'h3B3D] <= 28;
        weight_mem[16'h3B3E] <= 61;
        weight_mem[16'h3B3F] <= 35;
        weight_mem[16'h3B40] <= 29;
        weight_mem[16'h3B41] <= 2;
        weight_mem[16'h3B42] <= 246;
        weight_mem[16'h3B43] <= 248;
        weight_mem[16'h3B44] <= 253;
        weight_mem[16'h3B45] <= 21;
        weight_mem[16'h3B46] <= 39;
        weight_mem[16'h3B47] <= 32;
        weight_mem[16'h3B48] <= 35;
        weight_mem[16'h3B49] <= 61;
        weight_mem[16'h3B4A] <= 36;
        weight_mem[16'h3B4B] <= 37;
        weight_mem[16'h3B4C] <= 17;
        weight_mem[16'h3B4D] <= 238;
        weight_mem[16'h3B4E] <= 232;
        weight_mem[16'h3B4F] <= 253;
        weight_mem[16'h3B50] <= 238;
        weight_mem[16'h3B51] <= 243;
        weight_mem[16'h3B52] <= 235;
        weight_mem[16'h3B53] <= 248;
        weight_mem[16'h3B54] <= 240;
        weight_mem[16'h3B55] <= 3;
        weight_mem[16'h3B56] <= 241;
        weight_mem[16'h3B57] <= 242;
        weight_mem[16'h3B58] <= 7;
        weight_mem[16'h3B59] <= 24;
        weight_mem[16'h3B5A] <= 48;
        weight_mem[16'h3B5B] <= 45;
        weight_mem[16'h3B5C] <= 34;
        weight_mem[16'h3B5D] <= 34;
        weight_mem[16'h3B5E] <= 11;
        weight_mem[16'h3B5F] <= 13;
        weight_mem[16'h3B60] <= 26;
        weight_mem[16'h3B61] <= 31;
        weight_mem[16'h3B62] <= 21;
        weight_mem[16'h3B63] <= 22;
        weight_mem[16'h3B64] <= 241;
        weight_mem[16'h3B65] <= 252;
        weight_mem[16'h3B66] <= 247;
        weight_mem[16'h3B67] <= 253;
        weight_mem[16'h3B68] <= 235;
        weight_mem[16'h3B69] <= 248;
        weight_mem[16'h3B6A] <= 249;
        weight_mem[16'h3B6B] <= 242;
        weight_mem[16'h3B6C] <= 240;
        weight_mem[16'h3B6D] <= 237;
        weight_mem[16'h3B6E] <= 227;
        weight_mem[16'h3B6F] <= 248;
        weight_mem[16'h3B70] <= 2;
        weight_mem[16'h3B71] <= 18;
        weight_mem[16'h3B72] <= 29;
        weight_mem[16'h3B73] <= 48;
        weight_mem[16'h3B74] <= 27;
        weight_mem[16'h3B75] <= 30;
        weight_mem[16'h3B76] <= 7;
        weight_mem[16'h3B77] <= 248;
        weight_mem[16'h3B78] <= 243;
        weight_mem[16'h3B79] <= 1;
        weight_mem[16'h3B7A] <= 241;
        weight_mem[16'h3B7B] <= 249;
        weight_mem[16'h3B7C] <= 240;
        weight_mem[16'h3B7D] <= 252;
        weight_mem[16'h3B7E] <= 253;
        weight_mem[16'h3B7F] <= 237;
        weight_mem[16'h3B80] <= 247;
        weight_mem[16'h3B81] <= 237;
        weight_mem[16'h3B82] <= 234;
        weight_mem[16'h3B83] <= 245;
        weight_mem[16'h3B84] <= 227;
        weight_mem[16'h3B85] <= 226;
        weight_mem[16'h3B86] <= 245;
        weight_mem[16'h3B87] <= 227;
        weight_mem[16'h3B88] <= 244;
        weight_mem[16'h3B89] <= 248;
        weight_mem[16'h3B8A] <= 252;
        weight_mem[16'h3B8B] <= 0;
        weight_mem[16'h3B8C] <= 0;
        weight_mem[16'h3B8D] <= 245;
        weight_mem[16'h3B8E] <= 0;
        weight_mem[16'h3B8F] <= 245;
        weight_mem[16'h3B90] <= 244;
        weight_mem[16'h3B91] <= 247;
        weight_mem[16'h3B92] <= 232;
        weight_mem[16'h3B93] <= 253;
        weight_mem[16'h3B94] <= 247;
        weight_mem[16'h3B95] <= 249;
        weight_mem[16'h3B96] <= 232;
        weight_mem[16'h3B97] <= 247;
        weight_mem[16'h3B98] <= 237;
        weight_mem[16'h3B99] <= 235;
        weight_mem[16'h3B9A] <= 250;
        weight_mem[16'h3B9B] <= 241;
        weight_mem[16'h3B9C] <= 241;
        weight_mem[16'h3B9D] <= 236;
        weight_mem[16'h3B9E] <= 235;
        weight_mem[16'h3B9F] <= 231;
        weight_mem[16'h3BA0] <= 234;
        weight_mem[16'h3BA1] <= 239;
        weight_mem[16'h3BA2] <= 249;
        weight_mem[16'h3BA3] <= 241;
        weight_mem[16'h3BA4] <= 230;
        weight_mem[16'h3BA5] <= 241;
        weight_mem[16'h3BA6] <= 242;
        weight_mem[16'h3BA7] <= 241;
        weight_mem[16'h3BA8] <= 229;
        weight_mem[16'h3BA9] <= 240;
        weight_mem[16'h3BAA] <= 231;
        weight_mem[16'h3BAB] <= 230;
        weight_mem[16'h3BAC] <= 243;
        weight_mem[16'h3BAD] <= 233;
        weight_mem[16'h3BAE] <= 231;
        weight_mem[16'h3BAF] <= 235;

        // layer 2 neuron 0
        weight_mem[16'h4000] <= 11;
        weight_mem[16'h4001] <= 0;
        weight_mem[16'h4002] <= 5;
        weight_mem[16'h4003] <= 58;
        weight_mem[16'h4004] <= 3;
        weight_mem[16'h4005] <= 0;
        weight_mem[16'h4006] <= 79;
        weight_mem[16'h4007] <= 4;
        weight_mem[16'h4008] <= 247;
        weight_mem[16'h4009] <= 72;
        weight_mem[16'h400A] <= 0;
        weight_mem[16'h400B] <= 223;
        weight_mem[16'h400C] <= 247;
        weight_mem[16'h400D] <= 3;
        weight_mem[16'h400E] <= 5;
        weight_mem[16'h400F] <= 1;
        weight_mem[16'h4010] <= 5;
        weight_mem[16'h4011] <= 0;
        weight_mem[16'h4012] <= 3;
        weight_mem[16'h4013] <= 251;
        weight_mem[16'h4014] <= 0;
        weight_mem[16'h4015] <= 0;
        weight_mem[16'h4016] <= 0;
        weight_mem[16'h4017] <= 0;
        weight_mem[16'h4018] <= 127;
        weight_mem[16'h4019] <= 2;
        weight_mem[16'h401A] <= 14;
        weight_mem[16'h401B] <= 42;
        weight_mem[16'h401C] <= 2;
        weight_mem[16'h401D] <= 28;

        // layer 2 neuron 1
        weight_mem[16'h4200] <= 44;
        weight_mem[16'h4201] <= 0;
        weight_mem[16'h4202] <= 5;
        weight_mem[16'h4203] <= 225;
        weight_mem[16'h4204] <= 30;
        weight_mem[16'h4205] <= 0;
        weight_mem[16'h4206] <= 220;
        weight_mem[16'h4207] <= 4;
        weight_mem[16'h4208] <= 52;
        weight_mem[16'h4209] <= 37;
        weight_mem[16'h420A] <= 0;
        weight_mem[16'h420B] <= 51;
        weight_mem[16'h420C] <= 9;
        weight_mem[16'h420D] <= 251;
        weight_mem[16'h420E] <= 6;
        weight_mem[16'h420F] <= 253;
        weight_mem[16'h4210] <= 33;
        weight_mem[16'h4211] <= 0;
        weight_mem[16'h4212] <= 2;
        weight_mem[16'h4213] <= 208;
        weight_mem[16'h4214] <= 0;
        weight_mem[16'h4215] <= 3;
        weight_mem[16'h4216] <= 0;
        weight_mem[16'h4217] <= 0;
        weight_mem[16'h4218] <= 163;
        weight_mem[16'h4219] <= 211;
        weight_mem[16'h421A] <= 127;
        weight_mem[16'h421B] <= 238;
        weight_mem[16'h421C] <= 250;
        weight_mem[16'h421D] <= 12;

        // layer 2 neuron 2
        weight_mem[16'h4400] <= 174;
        weight_mem[16'h4401] <= 0;
        weight_mem[16'h4402] <= 252;
        weight_mem[16'h4403] <= 10;
        weight_mem[16'h4404] <= 21;
        weight_mem[16'h4405] <= 0;
        weight_mem[16'h4406] <= 25;
        weight_mem[16'h4407] <= 8;
        weight_mem[16'h4408] <= 9;
        weight_mem[16'h4409] <= 54;
        weight_mem[16'h440A] <= 0;
        weight_mem[16'h440B] <= 238;
        weight_mem[16'h440C] <= 5;
        weight_mem[16'h440D] <= 0;
        weight_mem[16'h440E] <= 2;
        weight_mem[16'h440F] <= 248;
        weight_mem[16'h4410] <= 81;
        weight_mem[16'h4411] <= 0;
        weight_mem[16'h4412] <= 255;
        weight_mem[16'h4413] <= 19;
        weight_mem[16'h4414] <= 0;
        weight_mem[16'h4415] <= 4;
        weight_mem[16'h4416] <= 0;
        weight_mem[16'h4417] <= 0;
        weight_mem[16'h4418] <= 204;
        weight_mem[16'h4419] <= 244;
        weight_mem[16'h441A] <= 235;
        weight_mem[16'h441B] <= 26;
        weight_mem[16'h441C] <= 255;
        weight_mem[16'h441D] <= 128;

        // layer 2 neuron 3
        weight_mem[16'h4600] <= 228;
        weight_mem[16'h4601] <= 0;
        weight_mem[16'h4602] <= 252;
        weight_mem[16'h4603] <= 243;
        weight_mem[16'h4604] <= 73;
        weight_mem[16'h4605] <= 0;
        weight_mem[16'h4606] <= 229;
        weight_mem[16'h4607] <= 247;
        weight_mem[16'h4608] <= 60;
        weight_mem[16'h4609] <= 128;
        weight_mem[16'h460A] <= 0;
        weight_mem[16'h460B] <= 69;
        weight_mem[16'h460C] <= 254;
        weight_mem[16'h460D] <= 6;
        weight_mem[16'h460E] <= 250;
        weight_mem[16'h460F] <= 255;
        weight_mem[16'h4610] <= 70;
        weight_mem[16'h4611] <= 0;
        weight_mem[16'h4612] <= 252;
        weight_mem[16'h4613] <= 54;
        weight_mem[16'h4614] <= 0;
        weight_mem[16'h4615] <= 252;
        weight_mem[16'h4616] <= 0;
        weight_mem[16'h4617] <= 0;
        weight_mem[16'h4618] <= 250;
        weight_mem[16'h4619] <= 79;
        weight_mem[16'h461A] <= 182;
        weight_mem[16'h461B] <= 229;
        weight_mem[16'h461C] <= 254;
        weight_mem[16'h461D] <= 44;

        // layer 2 neuron 4
        weight_mem[16'h4800] <= 61;
        weight_mem[16'h4801] <= 0;
        weight_mem[16'h4802] <= 6;
        weight_mem[16'h4803] <= 128;
        weight_mem[16'h4804] <= 252;
        weight_mem[16'h4805] <= 0;
        weight_mem[16'h4806] <= 196;
        weight_mem[16'h4807] <= 8;
        weight_mem[16'h4808] <= 22;
        weight_mem[16'h4809] <= 230;
        weight_mem[16'h480A] <= 0;
        weight_mem[16'h480B] <= 49;
        weight_mem[16'h480C] <= 1;
        weight_mem[16'h480D] <= 1;
        weight_mem[16'h480E] <= 6;
        weight_mem[16'h480F] <= 1;
        weight_mem[16'h4810] <= 1;
        weight_mem[16'h4811] <= 0;
        weight_mem[16'h4812] <= 252;
        weight_mem[16'h4813] <= 251;
        weight_mem[16'h4814] <= 0;
        weight_mem[16'h4815] <= 251;
        weight_mem[16'h4816] <= 0;
        weight_mem[16'h4817] <= 0;
        weight_mem[16'h4818] <= 225;
        weight_mem[16'h4819] <= 44;
        weight_mem[16'h481A] <= 74;
        weight_mem[16'h481B] <= 70;
        weight_mem[16'h481C] <= 0;
        weight_mem[16'h481D] <= 4;

        // layer 2 neuron 5
        weight_mem[16'h4A00] <= 0;
        weight_mem[16'h4A01] <= 0;
        weight_mem[16'h4A02] <= 0;
        weight_mem[16'h4A03] <= 0;
        weight_mem[16'h4A04] <= 0;
        weight_mem[16'h4A05] <= 0;
        weight_mem[16'h4A06] <= 254;
        weight_mem[16'h4A07] <= 0;
        weight_mem[16'h4A08] <= 129;
        weight_mem[16'h4A09] <= 254;
        weight_mem[16'h4A0A] <= 0;
        weight_mem[16'h4A0B] <= 0;
        weight_mem[16'h4A0C] <= 0;
        weight_mem[16'h4A0D] <= 0;
        weight_mem[16'h4A0E] <= 0;
        weight_mem[16'h4A0F] <= 0;
        weight_mem[16'h4A10] <= 241;
        weight_mem[16'h4A11] <= 0;
        weight_mem[16'h4A12] <= 0;
        weight_mem[16'h4A13] <= 0;
        weight_mem[16'h4A14] <= 0;
        weight_mem[16'h4A15] <= 0;
        weight_mem[16'h4A16] <= 0;
        weight_mem[16'h4A17] <= 0;
        weight_mem[16'h4A18] <= 0;
        weight_mem[16'h4A19] <= 0;
        weight_mem[16'h4A1A] <= 0;
        weight_mem[16'h4A1B] <= 0;
        weight_mem[16'h4A1C] <= 0;
        weight_mem[16'h4A1D] <= 0;

        // layer 2 neuron 6
        weight_mem[16'h4C00] <= 115;
        weight_mem[16'h4C01] <= 0;
        weight_mem[16'h4C02] <= 8;
        weight_mem[16'h4C03] <= 72;
        weight_mem[16'h4C04] <= 3;
        weight_mem[16'h4C05] <= 0;
        weight_mem[16'h4C06] <= 4;
        weight_mem[16'h4C07] <= 0;
        weight_mem[16'h4C08] <= 17;
        weight_mem[16'h4C09] <= 30;
        weight_mem[16'h4C0A] <= 0;
        weight_mem[16'h4C0B] <= 74;
        weight_mem[16'h4C0C] <= 5;
        weight_mem[16'h4C0D] <= 249;
        weight_mem[16'h4C0E] <= 4;
        weight_mem[16'h4C0F] <= 3;
        weight_mem[16'h4C10] <= 2;
        weight_mem[16'h4C11] <= 0;
        weight_mem[16'h4C12] <= 5;
        weight_mem[16'h4C13] <= 143;
        weight_mem[16'h4C14] <= 0;
        weight_mem[16'h4C15] <= 255;
        weight_mem[16'h4C16] <= 0;
        weight_mem[16'h4C17] <= 0;
        weight_mem[16'h4C18] <= 18;
        weight_mem[16'h4C19] <= 251;
        weight_mem[16'h4C1A] <= 108;
        weight_mem[16'h4C1B] <= 136;
        weight_mem[16'h4C1C] <= 252;
        weight_mem[16'h4C1D] <= 127;

        // layer 2 neuron 7
        weight_mem[16'h4E00] <= 63;
        weight_mem[16'h4E01] <= 0;
        weight_mem[16'h4E02] <= 1;
        weight_mem[16'h4E03] <= 117;
        weight_mem[16'h4E04] <= 149;
        weight_mem[16'h4E05] <= 0;
        weight_mem[16'h4E06] <= 240;
        weight_mem[16'h4E07] <= 255;
        weight_mem[16'h4E08] <= 25;
        weight_mem[16'h4E09] <= 14;
        weight_mem[16'h4E0A] <= 0;
        weight_mem[16'h4E0B] <= 223;
        weight_mem[16'h4E0C] <= 9;
        weight_mem[16'h4E0D] <= 249;
        weight_mem[16'h4E0E] <= 7;
        weight_mem[16'h4E0F] <= 5;
        weight_mem[16'h4E10] <= 88;
        weight_mem[16'h4E11] <= 0;
        weight_mem[16'h4E12] <= 4;
        weight_mem[16'h4E13] <= 27;
        weight_mem[16'h4E14] <= 0;
        weight_mem[16'h4E15] <= 4;
        weight_mem[16'h4E16] <= 0;
        weight_mem[16'h4E17] <= 0;
        weight_mem[16'h4E18] <= 158;
        weight_mem[16'h4E19] <= 27;
        weight_mem[16'h4E1A] <= 129;
        weight_mem[16'h4E1B] <= 59;
        weight_mem[16'h4E1C] <= 254;
        weight_mem[16'h4E1D] <= 7;

        // layer 2 neuron 8
        weight_mem[16'h5000] <= 211;
        weight_mem[16'h5001] <= 0;
        weight_mem[16'h5002] <= 255;
        weight_mem[16'h5003] <= 208;
        weight_mem[16'h5004] <= 128;
        weight_mem[16'h5005] <= 0;
        weight_mem[16'h5006] <= 39;
        weight_mem[16'h5007] <= 249;
        weight_mem[16'h5008] <= 83;
        weight_mem[16'h5009] <= 19;
        weight_mem[16'h500A] <= 0;
        weight_mem[16'h500B] <= 75;
        weight_mem[16'h500C] <= 12;
        weight_mem[16'h500D] <= 6;
        weight_mem[16'h500E] <= 255;
        weight_mem[16'h500F] <= 255;
        weight_mem[16'h5010] <= 39;
        weight_mem[16'h5011] <= 0;
        weight_mem[16'h5012] <= 251;
        weight_mem[16'h5013] <= 13;
        weight_mem[16'h5014] <= 0;
        weight_mem[16'h5015] <= 252;
        weight_mem[16'h5016] <= 0;
        weight_mem[16'h5017] <= 0;
        weight_mem[16'h5018] <= 98;
        weight_mem[16'h5019] <= 174;
        weight_mem[16'h501A] <= 224;
        weight_mem[16'h501B] <= 218;
        weight_mem[16'h501C] <= 249;
        weight_mem[16'h501D] <= 211;

        // layer 2 neuron 9
        weight_mem[16'h5200] <= 23;
        weight_mem[16'h5201] <= 0;
        weight_mem[16'h5202] <= 2;
        weight_mem[16'h5203] <= 17;
        weight_mem[16'h5204] <= 71;
        weight_mem[16'h5205] <= 0;
        weight_mem[16'h5206] <= 6;
        weight_mem[16'h5207] <= 9;
        weight_mem[16'h5208] <= 45;
        weight_mem[16'h5209] <= 65;
        weight_mem[16'h520A] <= 0;
        weight_mem[16'h520B] <= 10;
        weight_mem[16'h520C] <= 6;
        weight_mem[16'h520D] <= 251;
        weight_mem[16'h520E] <= 3;
        weight_mem[16'h520F] <= 0;
        weight_mem[16'h5210] <= 242;
        weight_mem[16'h5211] <= 0;
        weight_mem[16'h5212] <= 1;
        weight_mem[16'h5213] <= 175;
        weight_mem[16'h5214] <= 0;
        weight_mem[16'h5215] <= 1;
        weight_mem[16'h5216] <= 0;
        weight_mem[16'h5217] <= 0;
        weight_mem[16'h5218] <= 220;
        weight_mem[16'h5219] <= 222;
        weight_mem[16'h521A] <= 127;
        weight_mem[16'h521B] <= 211;
        weight_mem[16'h521C] <= 0;
        weight_mem[16'h521D] <= 193;

        // layer 2 neuron 10
        weight_mem[16'h5400] <= 215;
        weight_mem[16'h5401] <= 0;
        weight_mem[16'h5402] <= 245;
        weight_mem[16'h5403] <= 4;
        weight_mem[16'h5404] <= 127;
        weight_mem[16'h5405] <= 0;
        weight_mem[16'h5406] <= 69;
        weight_mem[16'h5407] <= 255;
        weight_mem[16'h5408] <= 80;
        weight_mem[16'h5409] <= 84;
        weight_mem[16'h540A] <= 0;
        weight_mem[16'h540B] <= 238;
        weight_mem[16'h540C] <= 251;
        weight_mem[16'h540D] <= 253;
        weight_mem[16'h540E] <= 0;
        weight_mem[16'h540F] <= 252;
        weight_mem[16'h5410] <= 244;
        weight_mem[16'h5411] <= 0;
        weight_mem[16'h5412] <= 0;
        weight_mem[16'h5413] <= 250;
        weight_mem[16'h5414] <= 0;
        weight_mem[16'h5415] <= 11;
        weight_mem[16'h5416] <= 0;
        weight_mem[16'h5417] <= 0;
        weight_mem[16'h5418] <= 184;
        weight_mem[16'h5419] <= 67;
        weight_mem[16'h541A] <= 43;
        weight_mem[16'h541B] <= 238;
        weight_mem[16'h541C] <= 0;
        weight_mem[16'h541D] <= 174;

        // layer 2 neuron 11
        weight_mem[16'h5600] <= 241;
        weight_mem[16'h5601] <= 0;
        weight_mem[16'h5602] <= 3;
        weight_mem[16'h5603] <= 240;
        weight_mem[16'h5604] <= 59;
        weight_mem[16'h5605] <= 0;
        weight_mem[16'h5606] <= 127;
        weight_mem[16'h5607] <= 2;
        weight_mem[16'h5608] <= 245;
        weight_mem[16'h5609] <= 227;
        weight_mem[16'h560A] <= 0;
        weight_mem[16'h560B] <= 232;
        weight_mem[16'h560C] <= 244;
        weight_mem[16'h560D] <= 4;
        weight_mem[16'h560E] <= 251;
        weight_mem[16'h560F] <= 5;
        weight_mem[16'h5610] <= 254;
        weight_mem[16'h5611] <= 0;
        weight_mem[16'h5612] <= 253;
        weight_mem[16'h5613] <= 57;
        weight_mem[16'h5614] <= 0;
        weight_mem[16'h5615] <= 8;
        weight_mem[16'h5616] <= 0;
        weight_mem[16'h5617] <= 0;
        weight_mem[16'h5618] <= 65;
        weight_mem[16'h5619] <= 75;
        weight_mem[16'h561A] <= 103;
        weight_mem[16'h561B] <= 213;
        weight_mem[16'h561C] <= 7;
        weight_mem[16'h561D] <= 19;

        // layer 2 neuron 12
        weight_mem[16'h5800] <= 58;
        weight_mem[16'h5801] <= 0;
        weight_mem[16'h5802] <= 1;
        weight_mem[16'h5803] <= 237;
        weight_mem[16'h5804] <= 205;
        weight_mem[16'h5805] <= 0;
        weight_mem[16'h5806] <= 23;
        weight_mem[16'h5807] <= 5;
        weight_mem[16'h5808] <= 42;
        weight_mem[16'h5809] <= 36;
        weight_mem[16'h580A] <= 0;
        weight_mem[16'h580B] <= 128;
        weight_mem[16'h580C] <= 6;
        weight_mem[16'h580D] <= 248;
        weight_mem[16'h580E] <= 12;
        weight_mem[16'h580F] <= 3;
        weight_mem[16'h5810] <= 27;
        weight_mem[16'h5811] <= 0;
        weight_mem[16'h5812] <= 3;
        weight_mem[16'h5813] <= 210;
        weight_mem[16'h5814] <= 0;
        weight_mem[16'h5815] <= 254;
        weight_mem[16'h5816] <= 0;
        weight_mem[16'h5817] <= 0;
        weight_mem[16'h5818] <= 169;
        weight_mem[16'h5819] <= 114;
        weight_mem[16'h581A] <= 149;
        weight_mem[16'h581B] <= 61;
        weight_mem[16'h581C] <= 254;
        weight_mem[16'h581D] <= 0;

        // layer 2 neuron 13
        weight_mem[16'h5A00] <= 242;
        weight_mem[16'h5A01] <= 0;
        weight_mem[16'h5A02] <= 240;
        weight_mem[16'h5A03] <= 43;
        weight_mem[16'h5A04] <= 127;
        weight_mem[16'h5A05] <= 0;
        weight_mem[16'h5A06] <= 230;
        weight_mem[16'h5A07] <= 254;
        weight_mem[16'h5A08] <= 35;
        weight_mem[16'h5A09] <= 47;
        weight_mem[16'h5A0A] <= 0;
        weight_mem[16'h5A0B] <= 60;
        weight_mem[16'h5A0C] <= 248;
        weight_mem[16'h5A0D] <= 1;
        weight_mem[16'h5A0E] <= 252;
        weight_mem[16'h5A0F] <= 244;
        weight_mem[16'h5A10] <= 6;
        weight_mem[16'h5A11] <= 0;
        weight_mem[16'h5A12] <= 1;
        weight_mem[16'h5A13] <= 9;
        weight_mem[16'h5A14] <= 0;
        weight_mem[16'h5A15] <= 249;
        weight_mem[16'h5A16] <= 0;
        weight_mem[16'h5A17] <= 0;
        weight_mem[16'h5A18] <= 58;
        weight_mem[16'h5A19] <= 248;
        weight_mem[16'h5A1A] <= 233;
        weight_mem[16'h5A1B] <= 79;
        weight_mem[16'h5A1C] <= 6;
        weight_mem[16'h5A1D] <= 198;

        // layer 2 neuron 14
        weight_mem[16'h5C00] <= 68;
        weight_mem[16'h5C01] <= 0;
        weight_mem[16'h5C02] <= 253;
        weight_mem[16'h5C03] <= 247;
        weight_mem[16'h5C04] <= 166;
        weight_mem[16'h5C05] <= 0;
        weight_mem[16'h5C06] <= 198;
        weight_mem[16'h5C07] <= 3;
        weight_mem[16'h5C08] <= 26;
        weight_mem[16'h5C09] <= 24;
        weight_mem[16'h5C0A] <= 0;
        weight_mem[16'h5C0B] <= 59;
        weight_mem[16'h5C0C] <= 250;
        weight_mem[16'h5C0D] <= 4;
        weight_mem[16'h5C0E] <= 2;
        weight_mem[16'h5C0F] <= 250;
        weight_mem[16'h5C10] <= 167;
        weight_mem[16'h5C11] <= 0;
        weight_mem[16'h5C12] <= 253;
        weight_mem[16'h5C13] <= 46;
        weight_mem[16'h5C14] <= 0;
        weight_mem[16'h5C15] <= 249;
        weight_mem[16'h5C16] <= 0;
        weight_mem[16'h5C17] <= 0;
        weight_mem[16'h5C18] <= 13;
        weight_mem[16'h5C19] <= 229;
        weight_mem[16'h5C1A] <= 207;
        weight_mem[16'h5C1B] <= 127;
        weight_mem[16'h5C1C] <= 7;
        weight_mem[16'h5C1D] <= 249;

        // layer 2 neuron 15
        weight_mem[16'h5E00] <= 228;
        weight_mem[16'h5E01] <= 0;
        weight_mem[16'h5E02] <= 255;
        weight_mem[16'h5E03] <= 5;
        weight_mem[16'h5E04] <= 110;
        weight_mem[16'h5E05] <= 0;
        weight_mem[16'h5E06] <= 238;
        weight_mem[16'h5E07] <= 248;
        weight_mem[16'h5E08] <= 25;
        weight_mem[16'h5E09] <= 192;
        weight_mem[16'h5E0A] <= 0;
        weight_mem[16'h5E0B] <= 170;
        weight_mem[16'h5E0C] <= 6;
        weight_mem[16'h5E0D] <= 254;
        weight_mem[16'h5E0E] <= 0;
        weight_mem[16'h5E0F] <= 3;
        weight_mem[16'h5E10] <= 80;
        weight_mem[16'h5E11] <= 0;
        weight_mem[16'h5E12] <= 255;
        weight_mem[16'h5E13] <= 222;
        weight_mem[16'h5E14] <= 0;
        weight_mem[16'h5E15] <= 3;
        weight_mem[16'h5E16] <= 0;
        weight_mem[16'h5E17] <= 0;
        weight_mem[16'h5E18] <= 128;
        weight_mem[16'h5E19] <= 48;
        weight_mem[16'h5E1A] <= 230;
        weight_mem[16'h5E1B] <= 238;
        weight_mem[16'h5E1C] <= 255;
        weight_mem[16'h5E1D] <= 108;

        // layer 3 neuron 0
        weight_mem[16'h8000] <= 78;
        weight_mem[16'h8001] <= 202;
        weight_mem[16'h8002] <= 57;
        weight_mem[16'h8003] <= 128;
        weight_mem[16'h8004] <= 183;
        weight_mem[16'h8005] <= 0;
        weight_mem[16'h8006] <= 187;
        weight_mem[16'h8007] <= 243;
        weight_mem[16'h8008] <= 227;
        weight_mem[16'h8009] <= 213;
        weight_mem[16'h800A] <= 193;
        weight_mem[16'h800B] <= 14;
        weight_mem[16'h800C] <= 188;
        weight_mem[16'h800D] <= 60;
        weight_mem[16'h800E] <= 70;
        weight_mem[16'h800F] <= 214;

        // layer 3 neuron 1
        weight_mem[16'h8200] <= 243;
        weight_mem[16'h8201] <= 75;
        weight_mem[16'h8202] <= 188;
        weight_mem[16'h8203] <= 42;
        weight_mem[16'h8204] <= 48;
        weight_mem[16'h8205] <= 0;
        weight_mem[16'h8206] <= 77;
        weight_mem[16'h8207] <= 136;
        weight_mem[16'h8208] <= 28;
        weight_mem[16'h8209] <= 37;
        weight_mem[16'h820A] <= 217;
        weight_mem[16'h820B] <= 15;
        weight_mem[16'h820C] <= 128;
        weight_mem[16'h820D] <= 176;
        weight_mem[16'h820E] <= 168;
        weight_mem[16'h820F] <= 39;

        // layer 3 neuron 2
        weight_mem[16'h8400] <= 254;
        weight_mem[16'h8401] <= 36;
        weight_mem[16'h8402] <= 18;
        weight_mem[16'h8403] <= 152;
        weight_mem[16'h8404] <= 78;
        weight_mem[16'h8405] <= 0;
        weight_mem[16'h8406] <= 28;
        weight_mem[16'h8407] <= 189;
        weight_mem[16'h8408] <= 20;
        weight_mem[16'h8409] <= 84;
        weight_mem[16'h840A] <= 29;
        weight_mem[16'h840B] <= 128;
        weight_mem[16'h840C] <= 38;
        weight_mem[16'h840D] <= 41;
        weight_mem[16'h840E] <= 35;
        weight_mem[16'h840F] <= 166;

        // layer 3 neuron 3
        weight_mem[16'h8600] <= 190;
        weight_mem[16'h8601] <= 17;
        weight_mem[16'h8602] <= 86;
        weight_mem[16'h8603] <= 233;
        weight_mem[16'h8604] <= 206;
        weight_mem[16'h8605] <= 0;
        weight_mem[16'h8606] <= 255;
        weight_mem[16'h8607] <= 184;
        weight_mem[16'h8608] <= 129;
        weight_mem[16'h8609] <= 86;
        weight_mem[16'h860A] <= 90;
        weight_mem[16'h860B] <= 4;
        weight_mem[16'h860C] <= 221;
        weight_mem[16'h860D] <= 52;
        weight_mem[16'h860E] <= 29;
        weight_mem[16'h860F] <= 46;

        // layer 3 neuron 4
        weight_mem[16'h8800] <= 219;
        weight_mem[16'h8801] <= 210;
        weight_mem[16'h8802] <= 128;
        weight_mem[16'h8803] <= 40;
        weight_mem[16'h8804] <= 44;
        weight_mem[16'h8805] <= 0;
        weight_mem[16'h8806] <= 198;
        weight_mem[16'h8807] <= 38;
        weight_mem[16'h8808] <= 190;
        weight_mem[16'h8809] <= 133;
        weight_mem[16'h880A] <= 220;
        weight_mem[16'h880B] <= 252;
        weight_mem[16'h880C] <= 74;
        weight_mem[16'h880D] <= 196;
        weight_mem[16'h880E] <= 26;
        weight_mem[16'h880F] <= 51;

        // layer 3 neuron 5
        weight_mem[16'h8A00] <= 4;
        weight_mem[16'h8A01] <= 128;
        weight_mem[16'h8A02] <= 246;
        weight_mem[16'h8A03] <= 70;
        weight_mem[16'h8A04] <= 224;
        weight_mem[16'h8A05] <= 0;
        weight_mem[16'h8A06] <= 182;
        weight_mem[16'h8A07] <= 190;
        weight_mem[16'h8A08] <= 21;
        weight_mem[16'h8A09] <= 216;
        weight_mem[16'h8A0A] <= 83;
        weight_mem[16'h8A0B] <= 70;
        weight_mem[16'h8A0C] <= 225;
        weight_mem[16'h8A0D] <= 32;
        weight_mem[16'h8A0E] <= 252;
        weight_mem[16'h8A0F] <= 239;

        // layer 3 neuron 6
        weight_mem[16'h8C00] <= 220;
        weight_mem[16'h8C01] <= 249;
        weight_mem[16'h8C02] <= 210;
        weight_mem[16'h8C03] <= 51;
        weight_mem[16'h8C04] <= 77;
        weight_mem[16'h8C05] <= 0;
        weight_mem[16'h8C06] <= 7;
        weight_mem[16'h8C07] <= 18;
        weight_mem[16'h8C08] <= 10;
        weight_mem[16'h8C09] <= 152;
        weight_mem[16'h8C0A] <= 128;
        weight_mem[16'h8C0B] <= 164;
        weight_mem[16'h8C0C] <= 212;
        weight_mem[16'h8C0D] <= 17;
        weight_mem[16'h8C0E] <= 65;
        weight_mem[16'h8C0F] <= 160;

        // layer 3 neuron 7
        weight_mem[16'h8E00] <= 69;
        weight_mem[16'h8E01] <= 75;
        weight_mem[16'h8E02] <= 148;
        weight_mem[16'h8E03] <= 128;
        weight_mem[16'h8E04] <= 13;
        weight_mem[16'h8E05] <= 0;
        weight_mem[16'h8E06] <= 80;
        weight_mem[16'h8E07] <= 32;
        weight_mem[16'h8E08] <= 224;
        weight_mem[16'h8E09] <= 24;
        weight_mem[16'h8E0A] <= 250;
        weight_mem[16'h8E0B] <= 65;
        weight_mem[16'h8E0C] <= 40;
        weight_mem[16'h8E0D] <= 156;
        weight_mem[16'h8E0E] <= 167;
        weight_mem[16'h8E0F] <= 200;

        // layer 3 neuron 8
        weight_mem[16'h9000] <= 178;
        weight_mem[16'h9001] <= 249;
        weight_mem[16'h9002] <= 121;
        weight_mem[16'h9003] <= 249;
        weight_mem[16'h9004] <= 242;
        weight_mem[16'h9005] <= 0;
        weight_mem[16'h9006] <= 175;
        weight_mem[16'h9007] <= 54;
        weight_mem[16'h9008] <= 65;
        weight_mem[16'h9009] <= 235;
        weight_mem[16'h900A] <= 32;
        weight_mem[16'h900B] <= 128;
        weight_mem[16'h900C] <= 35;
        weight_mem[16'h900D] <= 195;
        weight_mem[16'h900E] <= 221;
        weight_mem[16'h900F] <= 20;

        // layer 3 neuron 9
        weight_mem[16'h9200] <= 3;
        weight_mem[16'h9201] <= 218;
        weight_mem[16'h9202] <= 190;
        weight_mem[16'h9203] <= 9;
        weight_mem[16'h9204] <= 135;
        weight_mem[16'h9205] <= 0;
        weight_mem[16'h9206] <= 35;
        weight_mem[16'h9207] <= 52;
        weight_mem[16'h9208] <= 128;
        weight_mem[16'h9209] <= 216;
        weight_mem[16'h920A] <= 6;
        weight_mem[16'h920B] <= 191;
        weight_mem[16'h920C] <= 41;
        weight_mem[16'h920D] <= 1;
        weight_mem[16'h920E] <= 254;
        weight_mem[16'h920F] <= 97;
    end

    always @(posedge clk) begin
        if (reset) begin
            weight_val <= 0;
        end else begin 
            weight_val <= weight_mem[input_addr];
        end
    end

endmodule

