library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;entity weight_rom is    port(
        clk : in std_logic;
        totaladr: in unsigned(9 downto 0);
        weight : out signed(7 downto 0)
        );
end WeightRom;

architecture synth of WeightRom is
begin
    process (clk) begin
        if rising_edge(clk) then
            case totaladr is
                when "0000000000" => weight <= "00100110";
                when "0000000001" => weight <= "01101110";
                when "0000000010" => weight <= "00110000";
                when "0000000011" => weight <= "01011010";
                when "0000000100" => weight <= "01101001";
                when "0000000101" => weight <= "00000000";
                when "0000000110" => weight <= "01010101";
                when "0000000111" => weight <= "00000111";
                when "0000001000" => weight <= "00101000";
                when "0000001001" => weight <= "00001011";
                when "0000001010" => weight <= "00100100";
                when "0000001011" => weight <= "01011001";
                when "0000001100" => weight <= "00100011";
                when "0000001101" => weight <= "01110011";
                when "0000001110" => weight <= "01010000";
                when "0000001111" => weight <= "00110010";
                when "0000010000" => weight <= "00100101";
                when "0000010001" => weight <= "00110010";
                when "0000010010" => weight <= "01001111";
                when "0000010011" => weight <= "01110000";
                when "0000010100" => weight <= "00011111";
                when "0000010101" => weight <= "00001111";
                when "0000010110" => weight <= "00101110";
                when "0000010111" => weight <= "00110011";
                when "0000011000" => weight <= "01101111";
                when "0000011001" => weight <= "00000011";
                when "0000011010" => weight <= "00011000";
                when "0000011011" => weight <= "00101010";
                when "0000100000" => weight <= "01101110";
                when "0000100001" => weight <= "01100110";
                when "0000100010" => weight <= "01000100";
                when "0000100011" => weight <= "01011110";
                when "0000100100" => weight <= "00000101";
                when "0000100101" => weight <= "00100001";
                when "0000100110" => weight <= "01110111";
                when "0000100111" => weight <= "01111110";
                when "0000101000" => weight <= "00000100";
                when "0000101001" => weight <= "00111001";
                when "0000101010" => weight <= "01100001";
                when "0000101011" => weight <= "00101110";
                when "0000101100" => weight <= "01111010";
                when "0000101101" => weight <= "01101101";
                when "0000101110" => weight <= "01001110";
                when "0000101111" => weight <= "00101110";
                when "0000110000" => weight <= "01001110";
                when "0000110001" => weight <= "01110010";
                when "0000110010" => weight <= "00101101";
                when "0000110011" => weight <= "00110101";
                when "0000110100" => weight <= "01100010";
                when "0000110101" => weight <= "00010101";
                when "0000110110" => weight <= "00001101";
                when "0000110111" => weight <= "00001111";
                when "0000111000" => weight <= "00001111";
                when "0000111001" => weight <= "01010011";
                when "0000111010" => weight <= "00000110";
                when "0000111011" => weight <= "00000010";
                when "0001000000" => weight <= "01000101";
                when "0001000001" => weight <= "01110010";
                when "0001000010" => weight <= "00010110";
                when "0001000011" => weight <= "01111010";
                when "0001000100" => weight <= "00000101";
                when "0001000101" => weight <= "00001100";
                when "0001000110" => weight <= "01101101";
                when "0001000111" => weight <= "00101110";
                when "0001001000" => weight <= "00001001";
                when "0001001001" => weight <= "00001111";
                when "0001001010" => weight <= "00100111";
                when "0001001011" => weight <= "00001110";
                when "0001001100" => weight <= "01101110";
                when "0001001101" => weight <= "00110010";
                when "0001001110" => weight <= "01010100";
                when "0001001111" => weight <= "01011011";
                when "0001010000" => weight <= "01100000";
                when "0001010001" => weight <= "00010110";
                when "0001010010" => weight <= "01101100";
                when "0001010011" => weight <= "00011110";
                when "0001010100" => weight <= "01101001";
                when "0001010101" => weight <= "00011101";
                when "0001010110" => weight <= "01110100";
                when "0001010111" => weight <= "00101011";
                when "0001011000" => weight <= "01101100";
                when "0001011001" => weight <= "01111011";
                when "0001011010" => weight <= "01000101";
                when "0001011011" => weight <= "00010010";
                when "0001100000" => weight <= "01001100";
                when "0001100001" => weight <= "01010110";
                when "0001100010" => weight <= "01000010";
                when "0001100011" => weight <= "01101111";
                when "0001100100" => weight <= "00000111";
                when "0001100101" => weight <= "00010010";
                when "0001100110" => weight <= "01011101";
                when "0001100111" => weight <= "00111001";
                when "0001101000" => weight <= "00010100";
                when "0001101001" => weight <= "01011100";
                when "0001101010" => weight <= "01011011";
                when "0001101011" => weight <= "00001010";
                when "0001101100" => weight <= "01101100";
                when "0001101101" => weight <= "01000101";
                when "0001101110" => weight <= "01010001";
                when "0001101111" => weight <= "00100010";
                when "0001110000" => weight <= "10000000";
                when "0001110001" => weight <= "01011001";
                when "0001110010" => weight <= "01110110";
                when "0001110011" => weight <= "01100000";
                when "0001110100" => weight <= "00010010";
                when "0001110101" => weight <= "00000011";
                when "0001110110" => weight <= "01011010";
                when "0001110111" => weight <= "01001001";
                when "0001111000" => weight <= "00111011";
                when "0001111001" => weight <= "01110101";
                when "0001111010" => weight <= "00100011";
                when "0001111011" => weight <= "00000111";
                when "0010000000" => weight <= "00000110";
                when "0010000001" => weight <= "01101011";
                when "0010000010" => weight <= "01001001";
                when "0010000011" => weight <= "00111000";
                when "0010000100" => weight <= "00100011";
                when "0010000101" => weight <= "00001011";
                when "0010000110" => weight <= "00100101";
                when "0010000111" => weight <= "01001001";
                when "0010001000" => weight <= "00110010";
                when "0010001001" => weight <= "11111011";
                when "0010001010" => weight <= "01101110";
                when "0010001011" => weight <= "01000010";
                when "0010001100" => weight <= "00100001";
                when "0010001101" => weight <= "01100011";
                when "0010001110" => weight <= "01101000";
                when "0010001111" => weight <= "00111110";
                when "0010010000" => weight <= "01001100";
                when "0010010001" => weight <= "11111111";
                when "0010010010" => weight <= "00000100";
                when "0010010011" => weight <= "00010000";
                when "0010010100" => weight <= "00110110";
                when "0010010101" => weight <= "01101001";
                when "0010010110" => weight <= "00110000";
                when "0010010111" => weight <= "00001110";
                when "0010011000" => weight <= "01101101";
                when "0010011001" => weight <= "00101000";
                when "0010011010" => weight <= "01010010";
                when "0010011011" => weight <= "00100111";
                when "0010100000" => weight <= "00111110";
                when "0010100001" => weight <= "00100101";
                when "0010100010" => weight <= "00100011";
                when "0010100011" => weight <= "00100100";
                when "0010100100" => weight <= "01110101";
                when "0010100101" => weight <= "00100111";
                when "0010100110" => weight <= "01011110";
                when "0010100111" => weight <= "01000100";
                when "0010101000" => weight <= "01000111";
                when "0010101001" => weight <= "00011101";
                when "0010101010" => weight <= "01000010";
                when "0010101011" => weight <= "11100111";
                when "0010101100" => weight <= "11011101";
                when "0010101101" => weight <= "00011101";
                when "0010101110" => weight <= "00101111";
                when "0010101111" => weight <= "00010101";
                when "0010110000" => weight <= "11110110";
                when "0010110001" => weight <= "11101101";
                when "0010110010" => weight <= "11100110";
                when "0010110011" => weight <= "00110111";
                when "0010110100" => weight <= "11110000";
                when "0010110101" => weight <= "01010001";
                when "0010110110" => weight <= "00000100";
                when "0010110111" => weight <= "01000011";
                when "0010111000" => weight <= "00101011";
                when "0010111001" => weight <= "00110010";
                when "0010111010" => weight <= "00101101";
                when "0010111011" => weight <= "00110101";
                when "0011000000" => weight <= "01111011";
                when "0011000001" => weight <= "01010000";
                when "0011000010" => weight <= "01010000";
                when "0011000011" => weight <= "00011000";
                when "0011000100" => weight <= "00111110";
                when "0011000101" => weight <= "01001000";
                when "0011000110" => weight <= "01010011";
                when "0011000111" => weight <= "01010101";
                when "0011001000" => weight <= "01000011";
                when "0011001001" => weight <= "00001110";
                when "0011001010" => weight <= "11000000";
                when "0011001011" => weight <= "00001000";
                when "0011001100" => weight <= "10111110";
                when "0011001101" => weight <= "11010101";
                when "0011001110" => weight <= "11101110";
                when "0011001111" => weight <= "11010100";
                when "0011010000" => weight <= "11101010";
                when "0011010001" => weight <= "10011111";
                when "0011010010" => weight <= "00000111";
                when "0011010011" => weight <= "11110010";
                when "0011010100" => weight <= "11111011";
                when "0011010101" => weight <= "00101111";
                when "0011010110" => weight <= "00001011";
                when "0011010111" => weight <= "00001101";
                when "0011011000" => weight <= "00001111";
                when "0011011001" => weight <= "01100010";
                when "0011011010" => weight <= "01100110";
                when "0011011011" => weight <= "01001100";
                when "0011100000" => weight <= "01100010";
                when "0011100001" => weight <= "01110100";
                when "0011100010" => weight <= "00100101";
                when "0011100011" => weight <= "01000010";
                when "0011100100" => weight <= "00011010";
                when "0011100101" => weight <= "00011001";
                when "0011100110" => weight <= "01100000";
                when "0011100111" => weight <= "00000001";
                when "0011101000" => weight <= "00111000";
                when "0011101001" => weight <= "00110010";
                when "0011101010" => weight <= "00100000";
                when "0011101011" => weight <= "11101101";
                when "0011101100" => weight <= "11110101";
                when "0011101101" => weight <= "00001010";
                when "0011101110" => weight <= "00000010";
                when "0011101111" => weight <= "11010111";
                when "0011110000" => weight <= "11110001";
                when "0011110001" => weight <= "11101011";
                when "0011110010" => weight <= "10010011";
                when "0011110011" => weight <= "10101111";
                when "0011110100" => weight <= "10111001";
                when "0011110101" => weight <= "10111011";
                when "0011110110" => weight <= "01000111";
                when "0011110111" => weight <= "01010000";
                when "0011111000" => weight <= "01001100";
                when "0011111001" => weight <= "01111011";
                when "0011111010" => weight <= "01101011";
                when "0011111011" => weight <= "01010011";
                when "0100000000" => weight <= "00000111";
                when "0100000001" => weight <= "01000010";
                when "0100000010" => weight <= "00011101";
                when "0100000011" => weight <= "01011011";
                when "0100000100" => weight <= "00111011";
                when "0100000101" => weight <= "01100011";
                when "0100000110" => weight <= "01010011";
                when "0100000111" => weight <= "00000011";
                when "0100001000" => weight <= "11100001";
                when "0100001001" => weight <= "00001000";
                when "0100001010" => weight <= "00000001";
                when "0100001011" => weight <= "11100110";
                when "0100001100" => weight <= "11111101";
                when "0100001101" => weight <= "00010111";
                when "0100001110" => weight <= "11001101";
                when "0100001111" => weight <= "11100100";
                when "0100010000" => weight <= "11101001";
                when "0100010001" => weight <= "11110100";
                when "0100010010" => weight <= "11100011";
                when "0100010011" => weight <= "11100001";
                when "0100010100" => weight <= "11011100";
                when "0100010101" => weight <= "00000101";
                when "0100010110" => weight <= "00100001";
                when "0100010111" => weight <= "01011000";
                when "0100011000" => weight <= "00011001";
                when "0100011001" => weight <= "00010101";
                when "0100011010" => weight <= "00101110";
                when "0100011011" => weight <= "01011110";
                when "0100100000" => weight <= "01100000";
                when "0100100001" => weight <= "00101011";
                when "0100100010" => weight <= "00010011";
                when "0100100011" => weight <= "01011001";
                when "0100100100" => weight <= "00011011";
                when "0100100101" => weight <= "11111010";
                when "0100100110" => weight <= "11110110";
                when "0100100111" => weight <= "11100001";
                when "0100101000" => weight <= "00010001";
                when "0100101001" => weight <= "11110111";
                when "0100101010" => weight <= "11010010";
                when "0100101011" => weight <= "11011111";
                when "0100101100" => weight <= "11001011";
                when "0100101101" => weight <= "11111100";
                when "0100101110" => weight <= "00010101";
                when "0100101111" => weight <= "00010000";
                when "0100110000" => weight <= "11110110";
                when "0100110001" => weight <= "11100110";
                when "0100110010" => weight <= "10100000";
                when "0100110011" => weight <= "10011001";
                when "0100110100" => weight <= "11110111";
                when "0100110101" => weight <= "10111011";
                when "0100110110" => weight <= "10111000";
                when "0100110111" => weight <= "00011100";
                when "0100111000" => weight <= "00100110";
                when "0100111001" => weight <= "00100011";
                when "0100111010" => weight <= "01110100";
                when "0100111011" => weight <= "01110101";
                when "0101000000" => weight <= "00110011";
                when "0101000001" => weight <= "00101000";
                when "0101000010" => weight <= "00001000";
                when "0101000011" => weight <= "01110001";
                when "0101000100" => weight <= "00010110";
                when "0101000101" => weight <= "00011001";
                when "0101000110" => weight <= "00010100";
                when "0101000111" => weight <= "00100101";
                when "0101001000" => weight <= "10111111";
                when "0101001001" => weight <= "11011111";
                when "0101001010" => weight <= "11110000";
                when "0101001011" => weight <= "11011100";
                when "0101001100" => weight <= "00000000";
                when "0101001101" => weight <= "11011011";
                when "0101001110" => weight <= "00100010";
                when "0101001111" => weight <= "11111100";
                when "0101010000" => weight <= "11111110";
                when "0101010001" => weight <= "00010001";
                when "0101010010" => weight <= "00100000";
                when "0101010011" => weight <= "00000000";
                when "0101010100" => weight <= "10110010";
                when "0101010101" => weight <= "11010001";
                when "0101010110" => weight <= "11111011";
                when "0101010111" => weight <= "11111111";
                when "0101011000" => weight <= "11111101";
                when "0101011001" => weight <= "00110000";
                when "0101011010" => weight <= "00100110";
                when "0101011011" => weight <= "01100010";
                when "0101100000" => weight <= "00111000";
                when "0101100001" => weight <= "01000100";
                when "0101100010" => weight <= "00111011";
                when "0101100011" => weight <= "00010110";
                when "0101100100" => weight <= "01010100";
                when "0101100101" => weight <= "00010110";
                when "0101100110" => weight <= "11110110";
                when "0101100111" => weight <= "11100101";
                when "0101101000" => weight <= "10110110";
                when "0101101001" => weight <= "11000011";
                when "0101101010" => weight <= "00001011";
                when "0101101011" => weight <= "00001000";
                when "0101101100" => weight <= "00000011";
                when "0101101101" => weight <= "00011110";
                when "0101101110" => weight <= "00100001";
                when "0101101111" => weight <= "11110100";
                when "0101110000" => weight <= "00101000";
                when "0101110001" => weight <= "00011001";
                when "0101110010" => weight <= "00010110";
                when "0101110011" => weight <= "00001110";
                when "0101110100" => weight <= "11010110";
                when "0101110101" => weight <= "10111110";
                when "0101110110" => weight <= "10111110";
                when "0101110111" => weight <= "11011010";
                when "0101111000" => weight <= "00011010";
                when "0101111001" => weight <= "01011110";
                when "0101111010" => weight <= "01010110";
                when "0101111011" => weight <= "01100100";
                when "0110000000" => weight <= "01010000";
                when "0110000001" => weight <= "00011000";
                when "0110000010" => weight <= "01111010";
                when "0110000011" => weight <= "01100010";
                when "0110000100" => weight <= "01110101";
                when "0110000101" => weight <= "00011110";
                when "0110000110" => weight <= "11011010";
                when "0110000111" => weight <= "00011000";
                when "0110001000" => weight <= "00001101";
                when "0110001001" => weight <= "11101000";
                when "0110001010" => weight <= "00001101";
                when "0110001011" => weight <= "11100100";
                when "0110001100" => weight <= "11000010";
                when "0110001101" => weight <= "11110000";
                when "0110001110" => weight <= "01011101";
                when "0110001111" => weight <= "01000011";
                when "0110010000" => weight <= "00100100";
                when "0110010001" => weight <= "00110110";
                when "0110010010" => weight <= "11110011";
                when "0110010011" => weight <= "00010001";
                when "0110010100" => weight <= "11100001";
                when "0110010101" => weight <= "11111110";
                when "0110010110" => weight <= "10101000";
                when "0110010111" => weight <= "00010111";
                when "0110011000" => weight <= "01010010";
                when "0110011001" => weight <= "01100111";
                when "0110011010" => weight <= "00000011";
                when "0110011011" => weight <= "01010100";
                when "0110100000" => weight <= "01101000";
                when "0110100001" => weight <= "00000000";
                when "0110100010" => weight <= "00001000";
                when "0110100011" => weight <= "00001110";
                when "0110100100" => weight <= "01110111";
                when "0110100101" => weight <= "11100011";
                when "0110100110" => weight <= "11011100";
                when "0110100111" => weight <= "11100000";
                when "0110101000" => weight <= "10111000";
                when "0110101001" => weight <= "11111010";
                when "0110101010" => weight <= "00010110";
                when "0110101011" => weight <= "10111101";
                when "0110101100" => weight <= "00111111";
                when "0110101101" => weight <= "01011001";
                when "0110101110" => weight <= "00001101";
                when "0110101111" => weight <= "00110111";
                when "0110110000" => weight <= "00100000";
                when "0110110001" => weight <= "00010011";
                when "0110110010" => weight <= "11111111";
                when "0110110011" => weight <= "10111011";
                when "0110110100" => weight <= "00000000";
                when "0110110101" => weight <= "00000001";
                when "0110110110" => weight <= "10100010";
                when "0110110111" => weight <= "11001011";
                when "0110111000" => weight <= "00100000";
                when "0110111001" => weight <= "01100111";
                when "0110111010" => weight <= "00111011";
                when "0110111011" => weight <= "00110001";
                when "0111000000" => weight <= "01011001";
                when "0111000001" => weight <= "01110110";
                when "0111000010" => weight <= "00111011";
                when "0111000011" => weight <= "00001010";
                when "0111000100" => weight <= "00100100";
                when "0111000101" => weight <= "01001010";
                when "0111000110" => weight <= "11000100";
                when "0111000111" => weight <= "10111010";
                when "0111001000" => weight <= "11001001";
                when "0111001001" => weight <= "00010100";
                when "0111001010" => weight <= "11110011";
                when "0111001011" => weight <= "00110100";
                when "0111001100" => weight <= "11100011";
                when "0111001101" => weight <= "00010110";
                when "0111001110" => weight <= "00101111";
                when "0111001111" => weight <= "10011001";
                when "0111010000" => weight <= "01101010";
                when "0111010001" => weight <= "01001110";
                when "0111010010" => weight <= "11111101";
                when "0111010011" => weight <= "11100111";
                when "0111010100" => weight <= "11001001";
                when "0111010101" => weight <= "11110110";
                when "0111010110" => weight <= "10110010";
                when "0111010111" => weight <= "11111000";
                when "0111011000" => weight <= "01001000";
                when "0111011001" => weight <= "00011010";
                when "0111011010" => weight <= "00100101";
                when "0111011011" => weight <= "00111110";
                when "0111100000" => weight <= "01111010";
                when "0111100001" => weight <= "01010001";
                when "0111100010" => weight <= "01001100";
                when "0111100011" => weight <= "00010011";
                when "0111100100" => weight <= "00111101";
                when "0111100101" => weight <= "11101100";
                when "0111100110" => weight <= "11101111";
                when "0111100111" => weight <= "00000000";
                when "0111101000" => weight <= "10100000";
                when "0111101001" => weight <= "11110111";
                when "0111101010" => weight <= "11010111";
                when "0111101011" => weight <= "00101110";
                when "0111101100" => weight <= "01001011";
                when "0111101101" => weight <= "00011100";
                when "0111101110" => weight <= "01011111";
                when "0111101111" => weight <= "00111100";
                when "0111110000" => weight <= "01110000";
                when "0111110001" => weight <= "00001101";
                when "0111110010" => weight <= "11111101";
                when "0111110011" => weight <= "11110000";
                when "0111110100" => weight <= "11010000";
                when "0111110101" => weight <= "11101001";
                when "0111110110" => weight <= "00010001";
                when "0111110111" => weight <= "00010001";
                when "0111111000" => weight <= "11101101";
                when "0111111001" => weight <= "00000000";
                when "0111111010" => weight <= "00111000";
                when "0111111011" => weight <= "00111111";
                when "1000000000" => weight <= "00101111";
                when "1000000001" => weight <= "00111001";
                when "1000000010" => weight <= "01111011";
                when "1000000011" => weight <= "01100110";
                when "1000000100" => weight <= "01010101";
                when "1000000101" => weight <= "00100111";
                when "1000000110" => weight <= "11001010";
                when "1000000111" => weight <= "11100011";
                when "1000001000" => weight <= "11010001";
                when "1000001001" => weight <= "11110100";
                when "1000001010" => weight <= "11101111";
                when "1000001011" => weight <= "01000000";
                when "1000001100" => weight <= "00110100";
                when "1000001101" => weight <= "01111100";
                when "1000001110" => weight <= "01101101";
                when "1000001111" => weight <= "01000100";
                when "1000010000" => weight <= "00000100";
                when "1000010001" => weight <= "11011110";
                when "1000010010" => weight <= "11100110";
                when "1000010011" => weight <= "11000100";
                when "1000010100" => weight <= "11110000";
                when "1000010101" => weight <= "00000000";
                when "1000010110" => weight <= "11101100";
                when "1000010111" => weight <= "00010100";
                when "1000011000" => weight <= "01001010";
                when "1000011001" => weight <= "01001011";
                when "1000011010" => weight <= "01100101";
                when "1000011011" => weight <= "01001101";
                when "1000100000" => weight <= "01100011";
                when "1000100001" => weight <= "00110110";
                when "1000100010" => weight <= "00000100";
                when "1000100011" => weight <= "01011110";
                when "1000100100" => weight <= "11111110";
                when "1000100101" => weight <= "11110111";
                when "1000100110" => weight <= "11100101";
                when "1000100111" => weight <= "11110000";
                when "1000101000" => weight <= "10010001";
                when "1000101001" => weight <= "00011111";
                when "1000101010" => weight <= "11000110";
                when "1000101011" => weight <= "00001110";
                when "1000101100" => weight <= "01100001";
                when "1000101101" => weight <= "00000101";
                when "1000101110" => weight <= "00100100";
                when "1000101111" => weight <= "01011100";
                when "1000110000" => weight <= "00100011";
                when "1000110001" => weight <= "11011010";
                when "1000110010" => weight <= "11100101";
                when "1000110011" => weight <= "11000111";
                when "1000110100" => weight <= "11110001";
                when "1000110101" => weight <= "11001000";
                when "1000110110" => weight <= "00010110";
                when "1000110111" => weight <= "00010111";
                when "1000111000" => weight <= "11110111";
                when "1000111001" => weight <= "01111101";
                when "1000111010" => weight <= "01011100";
                when "1000111011" => weight <= "00011100";
                when "1001000000" => weight <= "00111111";
                when "1001000001" => weight <= "00010011";
                when "1001000010" => weight <= "01111100";
                when "1001000011" => weight <= "00010001";
                when "1001000100" => weight <= "01000100";
                when "1001000101" => weight <= "00000001";
                when "1001000110" => weight <= "10101001";
                when "1001000111" => weight <= "11100011";
                when "1001001000" => weight <= "11100001";
                when "1001001001" => weight <= "10101101";
                when "1001001010" => weight <= "00010001";
                when "1001001011" => weight <= "00000110";
                when "1001001100" => weight <= "00101100";
                when "1001001101" => weight <= "00000010";
                when "1001001110" => weight <= "00101101";
                when "1001001111" => weight <= "01010101";
                when "1001010000" => weight <= "00101110";
                when "1001010001" => weight <= "10111010";
                when "1001010010" => weight <= "11101111";
                when "1001010011" => weight <= "11001000";
                when "1001010100" => weight <= "00011011";
                when "1001010101" => weight <= "11011010";
                when "1001010110" => weight <= "00100100";
                when "1001010111" => weight <= "00100111";
                when "1001011000" => weight <= "00101101";
                when "1001011001" => weight <= "01110111";
                when "1001011010" => weight <= "01001110";
                when "1001011011" => weight <= "01111011";
                when "1001100000" => weight <= "00111000";
                when "1001100001" => weight <= "01010111";
                when "1001100010" => weight <= "00010111";
                when "1001100011" => weight <= "01100010";
                when "1001100100" => weight <= "00001101";
                when "1001100101" => weight <= "01000100";
                when "1001100110" => weight <= "11001011";
                when "1001100111" => weight <= "10101010";
                when "1001101000" => weight <= "11001100";
                when "1001101001" => weight <= "10111111";
                when "1001101010" => weight <= "11110100";
                when "1001101011" => weight <= "11110010";
                when "1001101100" => weight <= "11011101";
                when "1001101101" => weight <= "00101010";
                when "1001101110" => weight <= "11111000";
                when "1001101111" => weight <= "11010001";
                when "1001110000" => weight <= "11100100";
                when "1001110001" => weight <= "11001010";
                when "1001110010" => weight <= "11000011";
                when "1001110011" => weight <= "00010010";
                when "1001110100" => weight <= "00101100";
                when "1001110101" => weight <= "11100001";
                when "1001110110" => weight <= "00001011";
                when "1001110111" => weight <= "01001010";
                when "1001111000" => weight <= "00110110";
                when "1001111001" => weight <= "01000110";
                when "1001111010" => weight <= "00101101";
                when "1001111011" => weight <= "01001111";
                when "1010000000" => weight <= "01101111";
                when "1010000001" => weight <= "00011010";
                when "1010000010" => weight <= "00001110";
                when "1010000011" => weight <= "01110101";
                when "1010000100" => weight <= "01001101";
                when "1010000101" => weight <= "00100011";
                when "1010000110" => weight <= "11100110";
                when "1010000111" => weight <= "00010001";
                when "1010001000" => weight <= "11101011";
                when "1010001001" => weight <= "11110110";
                when "1010001010" => weight <= "11111000";
                when "1010001011" => weight <= "11000100";
                when "1010001100" => weight <= "11111111";
                when "1010001101" => weight <= "11001001";
                when "1010001110" => weight <= "00101000";
                when "1010001111" => weight <= "10111100";
                when "1010010000" => weight <= "11010111";
                when "1010010001" => weight <= "00010110";
                when "1010010010" => weight <= "00001100";
                when "1010010011" => weight <= "11110110";
                when "1010010100" => weight <= "00011111";
                when "1010010101" => weight <= "00010000";
                when "1010010110" => weight <= "11110011";
                when "1010010111" => weight <= "00001011";
                when "1010011000" => weight <= "01110011";
                when "1010011001" => weight <= "01001011";
                when "1010011010" => weight <= "00110000";
                when "1010011011" => weight <= "00011011";
                when "1010100000" => weight <= "00011010";
                when "1010100001" => weight <= "00011110";
                when "1010100010" => weight <= "00101001";
                when "1010100011" => weight <= "01111101";
                when "1010100100" => weight <= "00100100";
                when "1010100101" => weight <= "01000010";
                when "1010100110" => weight <= "11011000";
                when "1010100111" => weight <= "11001101";
                when "1010101000" => weight <= "11001101";
                when "1010101001" => weight <= "11000111";
                when "1010101010" => weight <= "11110110";
                when "1010101011" => weight <= "10100001";
                when "1010101100" => weight <= "11010100";
                when "1010101101" => weight <= "11001110";
                when "1010101110" => weight <= "11110000";
                when "1010101111" => weight <= "10111100";
                when "1010110000" => weight <= "11010010";
                when "1010110001" => weight <= "11011110";
                when "1010110010" => weight <= "00011100";
                when "1010110011" => weight <= "00010000";
                when "1010110100" => weight <= "00100000";
                when "1010110101" => weight <= "11111111";
                when "1010110110" => weight <= "00001100";
                when "1010110111" => weight <= "01100010";
                when "1010111000" => weight <= "00001010";
                when "1010111001" => weight <= "01001101";
                when "1010111010" => weight <= "01111001";
                when "1010111011" => weight <= "00010010";
                when "1011000000" => weight <= "01111110";
                when "1011000001" => weight <= "01110110";
                when "1011000010" => weight <= "01000010";
                when "1011000011" => weight <= "01101110";
                when "1011000100" => weight <= "01000110";
                when "1011000101" => weight <= "01010100";
                when "1011000110" => weight <= "00100001";
                when "1011000111" => weight <= "00110010";
                when "1011001000" => weight <= "00000010";
                when "1011001001" => weight <= "00001111";
                when "1011001010" => weight <= "00001001";
                when "1011001011" => weight <= "11101011";
                when "1011001100" => weight <= "11110011";
                when "1011001101" => weight <= "10111010";
                when "1011001110" => weight <= "10110100";
                when "1011001111" => weight <= "11110010";
                when "1011010000" => weight <= "00010001";
                when "1011010001" => weight <= "11010001";
                when "1011010010" => weight <= "11111000";
                when "1011010011" => weight <= "01000110";
                when "1011010100" => weight <= "11101011";
                when "1011010101" => weight <= "00010010";
                when "1011010110" => weight <= "00011000";
                when "1011010111" => weight <= "01001001";
                when "1011011000" => weight <= "00011010";
                when "1011011001" => weight <= "01101010";
                when "1011011010" => weight <= "01000110";
                when "1011011011" => weight <= "00100000";
                when "1011100000" => weight <= "00110000";
                when "1011100001" => weight <= "00000000";
                when "1011100010" => weight <= "00000010";
                when "1011100011" => weight <= "01010111";
                when "1011100100" => weight <= "01011011";
                when "1011100101" => weight <= "00110011";
                when "1011100110" => weight <= "01101010";
                when "1011100111" => weight <= "01000111";
                when "1011101000" => weight <= "00101111";
                when "1011101001" => weight <= "00110111";
                when "1011101010" => weight <= "00010010";
                when "1011101011" => weight <= "00000000";
                when "1011101100" => weight <= "10111010";
                when "1011101101" => weight <= "00000010";
                when "1011101110" => weight <= "11101100";
                when "1011101111" => weight <= "00101000";
                when "1011110000" => weight <= "00101110";
                when "1011110001" => weight <= "00011101";
                when "1011110010" => weight <= "01000010";
                when "1011110011" => weight <= "01001110";
                when "1011110100" => weight <= "01100001";
                when "1011110101" => weight <= "01100100";
                when "1011110110" => weight <= "00000000";
                when "1011110111" => weight <= "01101111";
                when "1011111000" => weight <= "00000010";
                when "1011111001" => weight <= "01100001";
                when "1011111010" => weight <= "01011010";
                when "1011111011" => weight <= "00010010";
                when "1100000000" => weight <= "00001000";
                when "1100000001" => weight <= "00010111";
                when "1100000010" => weight <= "00001010";
                when "1100000011" => weight <= "00110011";
                when "1100000100" => weight <= "01100100";
                when "1100000101" => weight <= "01011000";
                when "1100000110" => weight <= "01010011";
                when "1100000111" => weight <= "01110011";
                when "1100001000" => weight <= "01010110";
                when "1100001001" => weight <= "00101011";
                when "1100001010" => weight <= "00100001";
                when "1100001011" => weight <= "00101111";
                when "1100001100" => weight <= "01001000";
                when "1100001101" => weight <= "00100000";
                when "1100001110" => weight <= "01000010";
                when "1100001111" => weight <= "11111100";
                when "1100010000" => weight <= "01010001";
                when "1100010001" => weight <= "01011001";
                when "1100010010" => weight <= "01101100";
                when "1100010011" => weight <= "01011000";
                when "1100010100" => weight <= "01010110";
                when "1100010101" => weight <= "01100101";
                when "1100010110" => weight <= "00101101";
                when "1100010111" => weight <= "00001110";
                when "1100011000" => weight <= "00100001";
                when "1100011001" => weight <= "01100110";
                when "1100011010" => weight <= "01111100";
                when "1100011011" => weight <= "01000100";
                when "1100100000" => weight <= "00010011";
                when "1100100001" => weight <= "00000101";
                when "1100100010" => weight <= "01111011";
                when "1100100011" => weight <= "00010010";
                when "1100100100" => weight <= "01100011";
                when "1100100101" => weight <= "01110001";
                when "1100100110" => weight <= "01110101";
                when "1100100111" => weight <= "01001100";
                when "1100101000" => weight <= "01101100";
                when "1100101001" => weight <= "01101000";
                when "1100101010" => weight <= "01011011";
                when "1100101011" => weight <= "00101000";
                when "1100101100" => weight <= "01010100";
                when "1100101101" => weight <= "01100100";
                when "1100101110" => weight <= "00111101";
                when "1100101111" => weight <= "01001111";
                when "1100110000" => weight <= "01001110";
                when "1100110001" => weight <= "01001010";
                when "1100110010" => weight <= "01001110";
                when "1100110011" => weight <= "00101010";
                when "1100110100" => weight <= "01000100";
                when "1100110101" => weight <= "00111111";
                when "1100110110" => weight <= "00011001";
                when "1100110111" => weight <= "01101100";
                when "1100111000" => weight <= "00110110";
                when "1100111001" => weight <= "01010100";
                when "1100111010" => weight <= "01010110";
                when "1100111011" => weight <= "00100001";
                when "1101000000" => weight <= "00100010";
                when "1101000001" => weight <= "00100010";
                when "1101000010" => weight <= "01010010";
                when "1101000011" => weight <= "00110111";
                when "1101000100" => weight <= "01011001";
                when "1101000101" => weight <= "01100000";
                when "1101000110" => weight <= "00000111";
                when "1101000111" => weight <= "01100010";
                when "1101001000" => weight <= "01100110";
                when "1101001001" => weight <= "01001010";
                when "1101001010" => weight <= "00101000";
                when "1101001011" => weight <= "00111100";
                when "1101001100" => weight <= "01010000";
                when "1101001101" => weight <= "00110011";
                when "1101001110" => weight <= "01110011";
                when "1101001111" => weight <= "00011000";
                when "1101010000" => weight <= "01000011";
                when "1101010001" => weight <= "00010100";
                when "1101010010" => weight <= "00111101";
                when "1101010011" => weight <= "00101010";
                when "1101010100" => weight <= "00011111";
                when "1101010101" => weight <= "01000001";
                when "1101010110" => weight <= "01011101";
                when "1101010111" => weight <= "01011101";
                when "1101011000" => weight <= "00101001";
                when "1101011001" => weight <= "01001001";
                when "1101011010" => weight <= "01001001";
                when "1101011011" => weight <= "01100010";
                when "1101100000" => weight <= "00010011";
                when "1101100001" => weight <= "00111000";
                when "1101100010" => weight <= "01011101";
                when "1101100011" => weight <= "00100000";
                when "1101100100" => weight <= "00001011";
                when "1101100101" => weight <= "01101010";
                when "1101100110" => weight <= "01111110";
                when "1101100111" => weight <= "01110011";
                when "1101101000" => weight <= "01001101";
                when "1101101001" => weight <= "00010001";
                when "1101101010" => weight <= "00010110";
                when "1101101011" => weight <= "00100010";
                when "1101101100" => weight <= "00011101";
                when "1101101101" => weight <= "00011000";
                when "1101101110" => weight <= "01000101";
                when "1101101111" => weight <= "00000101";
                when "1101110000" => weight <= "01001110";
                when "1101110001" => weight <= "00000000";
                when "1101110010" => weight <= "01110011";
                when "1101110011" => weight <= "00100011";
                when "1101110100" => weight <= "01101010";
                when "1101110101" => weight <= "00100111";
                when "1101110110" => weight <= "00110000";
                when "1101110111" => weight <= "00111000";
                when "1101111000" => weight <= "01000000";
                when "1101111001" => weight <= "01011111";
                when "1101111010" => weight <= "00011110";
                when "1101111011" => weight <= "00010011";
                when others => weight <= "00000000";
        end case;
    end if;
    end process;
end;
