library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity digits_rom is
    Port ( address : in  STD_LOGIC_VECTOR(7 downto 0);
           data : out STD_LOGIC_VECTOR(5 downto 0));
end rom;

architecture Behavioral of rom is
begin
    process(address)
    begin
        case address is
            when "00000000" => data <= "111111";
            when "00000001" => data <= "111111";
            when "00000010" => data <= "111111";
            when "00000011" => data <= "000000";
            when "00000100" => data <= "000000";
            when "00000101" => data <= "111111";
            when "00000110" => data <= "000000";
            when "00000111" => data <= "000000";
            when "00001000" => data <= "111111";
            when "00001001" => data <= "111111";
            when "00001010" => data <= "111111";
            when "00001011" => data <= "000000";
            when "00001100" => data <= "111111";
            when "00001101" => data <= "111111";
            when "00001110" => data <= "111111";
            when "00001111" => data <= "000000";
            when "00010000" => data <= "111111";
            when "00010001" => data <= "000000";
            when "00010010" => data <= "000000";
            when "00010011" => data <= "000000";
            when "00010100" => data <= "111111";
            when "00010101" => data <= "111111";
            when "00010110" => data <= "111111";
            when "00010111" => data <= "000000";
            when "00011000" => data <= "111111";
            when "00011001" => data <= "000000";
            when "00011010" => data <= "000000";
            when "00011011" => data <= "000000";
            when "00011100" => data <= "111111";
            when "00011101" => data <= "111111";
            when "00011110" => data <= "111111";
            when "00011111" => data <= "000000";
            when "00100000" => data <= "111111";
            when "00100001" => data <= "111111";
            when "00100010" => data <= "111111";
            when "00100011" => data <= "000000";
            when "00100100" => data <= "111111";
            when "00100101" => data <= "111111";
            when "00100110" => data <= "111111";
            when "00100111" => data <= "000000";
            when "01000000" => data <= "111111";
            when "01000001" => data <= "000000";
            when "01000010" => data <= "111111";
            when "01000011" => data <= "000000";
            when "01000100" => data <= "111111";
            when "01000101" => data <= "111111";
            when "01000110" => data <= "000000";
            when "01000111" => data <= "000000";
            when "01001000" => data <= "000000";
            when "01001001" => data <= "000000";
            when "01001010" => data <= "111111";
            when "01001011" => data <= "000000";
            when "01001100" => data <= "000000";
            when "01001101" => data <= "111111";
            when "01001110" => data <= "111111";
            when "01001111" => data <= "000000";
            when "01010000" => data <= "111111";
            when "01010001" => data <= "000000";
            when "01010010" => data <= "111111";
            when "01010011" => data <= "000000";
            when "01010100" => data <= "111111";
            when "01010101" => data <= "000000";
            when "01010110" => data <= "000000";
            when "01010111" => data <= "000000";
            when "01011000" => data <= "111111";
            when "01011001" => data <= "111111";
            when "01011010" => data <= "111111";
            when "01011011" => data <= "000000";
            when "01011100" => data <= "000000";
            when "01011101" => data <= "000000";
            when "01011110" => data <= "111111";
            when "01011111" => data <= "000000";
            when "01100000" => data <= "111111";
            when "01100001" => data <= "000000";
            when "01100010" => data <= "111111";
            when "01100011" => data <= "000000";
            when "01100100" => data <= "111111";
            when "01100101" => data <= "000000";
            when "01100110" => data <= "111111";
            when "01100111" => data <= "000000";
            when "10000000" => data <= "111111";
            when "10000001" => data <= "000000";
            when "10000010" => data <= "111111";
            when "10000011" => data <= "000000";
            when "10000100" => data <= "000000";
            when "10000101" => data <= "111111";
            when "10000110" => data <= "000000";
            when "10000111" => data <= "000000";
            when "10001000" => data <= "111111";
            when "10001001" => data <= "111111";
            when "10001010" => data <= "000000";
            when "10001011" => data <= "000000";
            when "10001100" => data <= "000000";
            when "10001101" => data <= "000000";
            when "10001110" => data <= "111111";
            when "10001111" => data <= "000000";
            when "10010000" => data <= "111111";
            when "10010001" => data <= "111111";
            when "10010010" => data <= "111111";
            when "10010011" => data <= "000000";
            when "10010100" => data <= "000000";
            when "10010101" => data <= "111111";
            when "10010110" => data <= "111111";
            when "10010111" => data <= "000000";
            when "10011000" => data <= "111111";
            when "10011001" => data <= "000000";
            when "10011010" => data <= "111111";
            when "10011011" => data <= "000000";
            when "10011100" => data <= "000000";
            when "10011101" => data <= "000000";
            when "10011110" => data <= "111111";
            when "10011111" => data <= "000000";
            when "10100000" => data <= "111111";
            when "10100001" => data <= "111111";
            when "10100010" => data <= "111111";
            when "10100011" => data <= "000000";
            when "10100100" => data <= "111111";
            when "10100101" => data <= "111111";
            when "10100110" => data <= "111111";
            when "10100111" => data <= "000000";
            when "11000000" => data <= "111111";
            when "11000001" => data <= "111111";
            when "11000010" => data <= "111111";
            when "11000011" => data <= "000000";
            when "11000100" => data <= "000000";
            when "11000101" => data <= "111111";
            when "11000110" => data <= "000000";
            when "11000111" => data <= "000000";
            when "11001000" => data <= "111111";
            when "11001001" => data <= "111111";
            when "11001010" => data <= "111111";
            when "11001011" => data <= "000000";
            when "11001100" => data <= "111111";
            when "11001101" => data <= "111111";
            when "11001110" => data <= "111111";
            when "11001111" => data <= "000000";
            when "11010000" => data <= "000000";
            when "11010001" => data <= "000000";
            when "11010010" => data <= "111111";
            when "11010011" => data <= "000000";
            when "11010100" => data <= "111111";
            when "11010101" => data <= "111111";
            when "11010110" => data <= "111111";
            when "11010111" => data <= "000000";
            when "11011000" => data <= "111111";
            when "11011001" => data <= "111111";
            when "11011010" => data <= "111111";
            when "11011011" => data <= "000000";
            when "11011100" => data <= "000000";
            when "11011101" => data <= "000000";
            when "11011110" => data <= "111111";
            when "11011111" => data <= "000000";
            when "11100000" => data <= "111111";
            when "11100001" => data <= "111111";
            when "11100010" => data <= "111111";
            when "11100011" => data <= "000000";
            when "11100100" => data <= "000000";
            when "11100101" => data <= "000000";
            when "11100110" => data <= "111111";
            when "11100111" => data <= "000000";
            when others => data <= "000000";
        end case;
    end process;
end Behavioral;