library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;entity im3_1 is    port(
        clk : in std_logic;
        totaladr: in unsigned(3 downto 0);
        grayScale : out std_logic_vector(7 downto 0)
        );
end im3_1;

architecture synth of im3_1 is
begin
    process (clk) begin
        if rising_edge(clk) then
            case totaladr is
                when "0000" => grayScale <= "00000000";
                when "0001" => grayScale <= "00000000";
                when "0010" => grayScale <= "00000000";
                when "0011" => grayScale <= "00000000";
                when "00100" => grayScale <= "00000000";
                when "00101" => grayScale <= "00000000";
                when "00110" => grayScale <= "00000000";
                when "00111" => grayScale <= "00000000";
                when "001000" => grayScale <= "00000000";
                when "001001" => grayScale <= "00000000";
                when "001010" => grayScale <= "00000000";
                when "001011" => grayScale <= "00000000";
                when "001100" => grayScale <= "00000000";
                when "001101" => grayScale <= "00000000";
                when "001110" => grayScale <= "00000000";
                when "001111" => grayScale <= "00000000";
                when "0010000" => grayScale <= "00000000";
                when "0010001" => grayScale <= "00000000";
                when "0010010" => grayScale <= "00000000";
                when "0010011" => grayScale <= "00000000";
                when "0010100" => grayScale <= "00000000";
                when "0010101" => grayScale <= "00000000";
                when "0010110" => grayScale <= "00000000";
                when "0010111" => grayScale <= "00000000";
                when "0011000" => grayScale <= "00000000";
                when "0011001" => grayScale <= "00000000";
                when "0011010" => grayScale <= "00000000";
                when "0011011" => grayScale <= "00000000";
                when "0100" => grayScale <= "00000000";
                when "0101" => grayScale <= "00000000";
                when "0110" => grayScale <= "00000000";
                when "0111" => grayScale <= "00000000";
                when "01100" => grayScale <= "00000000";
                when "01101" => grayScale <= "00000000";
                when "01110" => grayScale <= "00000000";
                when "01111" => grayScale <= "00000000";
                when "011000" => grayScale <= "00000000";
                when "011001" => grayScale <= "00000000";
                when "011010" => grayScale <= "00000000";
                when "011011" => grayScale <= "00000000";
                when "011100" => grayScale <= "00000000";
                when "011101" => grayScale <= "00000000";
                when "011110" => grayScale <= "00000000";
                when "011111" => grayScale <= "00000000";
                when "0110000" => grayScale <= "00000000";
                when "0110001" => grayScale <= "00000000";
                when "0110010" => grayScale <= "00000000";
                when "0110011" => grayScale <= "00000000";
                when "0110100" => grayScale <= "00000000";
                when "0110101" => grayScale <= "00000000";
                when "0110110" => grayScale <= "00000000";
                when "0110111" => grayScale <= "00000000";
                when "0111000" => grayScale <= "00000000";
                when "0111001" => grayScale <= "00000000";
                when "0111010" => grayScale <= "00000000";
                when "0111011" => grayScale <= "00000000";
                when "1000" => grayScale <= "00000000";
                when "1001" => grayScale <= "00000000";
                when "1010" => grayScale <= "00000000";
                when "1011" => grayScale <= "00000000";
                when "10100" => grayScale <= "00000000";
                when "10101" => grayScale <= "00000000";
                when "10110" => grayScale <= "00000000";
                when "10111" => grayScale <= "00000000";
                when "101000" => grayScale <= "00000000";
                when "101001" => grayScale <= "00000000";
                when "101010" => grayScale <= "00000000";
                when "101011" => grayScale <= "00000000";
                when "101100" => grayScale <= "00000000";
                when "101101" => grayScale <= "00000000";
                when "101110" => grayScale <= "00000000";
                when "101111" => grayScale <= "00000000";
                when "1010000" => grayScale <= "00000000";
                when "1010001" => grayScale <= "00000000";
                when "1010010" => grayScale <= "00000000";
                when "1010011" => grayScale <= "00000000";
                when "1010100" => grayScale <= "00000000";
                when "1010101" => grayScale <= "00000000";
                when "1010110" => grayScale <= "00000000";
                when "1010111" => grayScale <= "00000000";
                when "1011000" => grayScale <= "00000000";
                when "1011001" => grayScale <= "00000000";
                when "1011010" => grayScale <= "00000000";
                when "1011011" => grayScale <= "00000000";
                when "1100" => grayScale <= "00000000";
                when "1101" => grayScale <= "00000000";
                when "1110" => grayScale <= "00000000";
                when "1111" => grayScale <= "00000000";
                when "11100" => grayScale <= "00000000";
                when "11101" => grayScale <= "00000000";
                when "11110" => grayScale <= "00000000";
                when "11111" => grayScale <= "00000000";
                when "111000" => grayScale <= "00000000";
                when "111001" => grayScale <= "00000000";
                when "111010" => grayScale <= "00000000";
                when "111011" => grayScale <= "00000000";
                when "111100" => grayScale <= "00000000";
                when "111101" => grayScale <= "00000000";
                when "111110" => grayScale <= "00000000";
                when "111111" => grayScale <= "00000000";
                when "1110000" => grayScale <= "00000000";
                when "1110001" => grayScale <= "00000000";
                when "1110010" => grayScale <= "00000000";
                when "1110011" => grayScale <= "00000000";
                when "1110100" => grayScale <= "00000000";
                when "1110101" => grayScale <= "00000000";
                when "1110110" => grayScale <= "00000000";
                when "1110111" => grayScale <= "00000000";
                when "1111000" => grayScale <= "00000000";
                when "1111001" => grayScale <= "00000000";
                when "1111010" => grayScale <= "00000000";
                when "1111011" => grayScale <= "00000000";
                when "10000" => grayScale <= "00000000";
                when "10001" => grayScale <= "00000000";
                when "10010" => grayScale <= "00000000";
                when "10011" => grayScale <= "00000000";
                when "100100" => grayScale <= "00000000";
                when "100101" => grayScale <= "00000000";
                when "100110" => grayScale <= "00000000";
                when "100111" => grayScale <= "00000000";
                when "1001000" => grayScale <= "00000000";
                when "1001001" => grayScale <= "00000000";
                when "1001010" => grayScale <= "00000000";
                when "1001011" => grayScale <= "00000000";
                when "1001100" => grayScale <= "00000000";
                when "1001101" => grayScale <= "00000000";
                when "1001110" => grayScale <= "00000000";
                when "1001111" => grayScale <= "00000000";
                when "10010000" => grayScale <= "00000000";
                when "10010001" => grayScale <= "00000000";
                when "10010010" => grayScale <= "01101101";
                when "10010011" => grayScale <= "01111110";
                when "10010100" => grayScale <= "01010101";
                when "10010101" => grayScale <= "00000000";
                when "10010110" => grayScale <= "00000000";
                when "10010111" => grayScale <= "00000000";
                when "10011000" => grayScale <= "00000000";
                when "10011001" => grayScale <= "00000000";
                when "10011010" => grayScale <= "00000000";
                when "10011011" => grayScale <= "00000000";
                when "10100" => grayScale <= "00000000";
                when "10101" => grayScale <= "00000000";
                when "10110" => grayScale <= "00000000";
                when "10111" => grayScale <= "00000000";
                when "101100" => grayScale <= "00000000";
                when "101101" => grayScale <= "00000000";
                when "101110" => grayScale <= "00000000";
                when "101111" => grayScale <= "00000000";
                when "1011000" => grayScale <= "00000000";
                when "1011001" => grayScale <= "00000000";
                when "1011010" => grayScale <= "00000000";
                when "1011011" => grayScale <= "00000000";
                when "1011100" => grayScale <= "00000000";
                when "1011101" => grayScale <= "00000000";
                when "1011110" => grayScale <= "00000000";
                when "1011111" => grayScale <= "00000000";
                when "10110000" => grayScale <= "00000000";
                when "10110001" => grayScale <= "00101111";
                when "10110010" => grayScale <= "01111011";
                when "10110011" => grayScale <= "01111110";
                when "10110100" => grayScale <= "01111110";
                when "10110101" => grayScale <= "00000000";
                when "10110110" => grayScale <= "00000000";
                when "10110111" => grayScale <= "00000000";
                when "10111000" => grayScale <= "00000000";
                when "10111001" => grayScale <= "00000000";
                when "10111010" => grayScale <= "00000000";
                when "10111011" => grayScale <= "00000000";
                when "11000" => grayScale <= "00000000";
                when "11001" => grayScale <= "00000000";
                when "11010" => grayScale <= "00000000";
                when "11011" => grayScale <= "00000000";
                when "110100" => grayScale <= "00000000";
                when "110101" => grayScale <= "00000000";
                when "110110" => grayScale <= "00000000";
                when "110111" => grayScale <= "00000000";
                when "1101000" => grayScale <= "00000000";
                when "1101001" => grayScale <= "00000000";
                when "1101010" => grayScale <= "00000000";
                when "1101011" => grayScale <= "00000000";
                when "1101100" => grayScale <= "00000000";
                when "1101101" => grayScale <= "00000000";
                when "1101110" => grayScale <= "00000000";
                when "1101111" => grayScale <= "00000000";
                when "11010000" => grayScale <= "00001010";
                when "11010001" => grayScale <= "01101010";
                when "11010010" => grayScale <= "01111110";
                when "11010011" => grayScale <= "01111011";
                when "11010100" => grayScale <= "01000010";
                when "11010101" => grayScale <= "00000000";
                when "11010110" => grayScale <= "00000000";
                when "11010111" => grayScale <= "00000000";
                when "11011000" => grayScale <= "00000000";
                when "11011001" => grayScale <= "00000000";
                when "11011010" => grayScale <= "00000000";
                when "11011011" => grayScale <= "00000000";
                when "11100" => grayScale <= "00000000";
                when "11101" => grayScale <= "00000000";
                when "11110" => grayScale <= "00000000";
                when "11111" => grayScale <= "00000000";
                when "111100" => grayScale <= "00000000";
                when "111101" => grayScale <= "00000000";
                when "111110" => grayScale <= "00000000";
                when "111111" => grayScale <= "00000000";
                when "1111000" => grayScale <= "00000000";
                when "1111001" => grayScale <= "00000000";
                when "1111010" => grayScale <= "00000000";
                when "1111011" => grayScale <= "00000000";
                when "1111100" => grayScale <= "00000000";
                when "1111101" => grayScale <= "00000000";
                when "1111110" => grayScale <= "00000000";
                when "1111111" => grayScale <= "00000000";
                when "11110000" => grayScale <= "01001000";
                when "11110001" => grayScale <= "01111110";
                when "11110010" => grayScale <= "01111110";
                when "11110011" => grayScale <= "01101011";
                when "11110100" => grayScale <= "00000000";
                when "11110101" => grayScale <= "00000000";
                when "11110110" => grayScale <= "00000000";
                when "11110111" => grayScale <= "00000000";
                when "11111000" => grayScale <= "00000000";
                when "11111001" => grayScale <= "00000000";
                when "11111010" => grayScale <= "00000000";
                when "11111011" => grayScale <= "00000000";
                when "100000" => grayScale <= "00000000";
                when "100001" => grayScale <= "00000000";
                when "100010" => grayScale <= "00000000";
                when "100011" => grayScale <= "00000000";
                when "1000100" => grayScale <= "00000000";
                when "1000101" => grayScale <= "00000000";
                when "1000110" => grayScale <= "00000000";
                when "1000111" => grayScale <= "00000000";
                when "10001000" => grayScale <= "00000000";
                when "10001001" => grayScale <= "00000000";
                when "10001010" => grayScale <= "00000000";
                when "10001011" => grayScale <= "00000000";
                when "10001100" => grayScale <= "00000000";
                when "10001101" => grayScale <= "00000000";
                when "10001110" => grayScale <= "00000000";
                when "10001111" => grayScale <= "00001000";
                when "100010000" => grayScale <= "01011111";
                when "100010001" => grayScale <= "01111110";
                when "100010010" => grayScale <= "01111110";
                when "100010011" => grayScale <= "01001100";
                when "100010100" => grayScale <= "00000000";
                when "100010101" => grayScale <= "00000000";
                when "100010110" => grayScale <= "00000000";
                when "100010111" => grayScale <= "00000000";
                when "100011000" => grayScale <= "00000000";
                when "100011001" => grayScale <= "00000000";
                when "100011010" => grayScale <= "00000000";
                when "100011011" => grayScale <= "00000000";
                when "100100" => grayScale <= "00000000";
                when "100101" => grayScale <= "00000000";
                when "100110" => grayScale <= "00000000";
                when "100111" => grayScale <= "00000000";
                when "1001100" => grayScale <= "00000000";
                when "1001101" => grayScale <= "00000000";
                when "1001110" => grayScale <= "00000000";
                when "1001111" => grayScale <= "00000000";
                when "10011000" => grayScale <= "00000000";
                when "10011001" => grayScale <= "00000000";
                when "10011010" => grayScale <= "00000000";
                when "10011011" => grayScale <= "00000000";
                when "10011100" => grayScale <= "00000000";
                when "10011101" => grayScale <= "00000000";
                when "10011110" => grayScale <= "00001010";
                when "10011111" => grayScale <= "01011010";
                when "100110000" => grayScale <= "01111110";
                when "100110001" => grayScale <= "01111110";
                when "100110010" => grayScale <= "01110011";
                when "100110011" => grayScale <= "00011001";
                when "100110100" => grayScale <= "00000000";
                when "100110101" => grayScale <= "00000000";
                when "100110110" => grayScale <= "00000000";
                when "100110111" => grayScale <= "00000000";
                when "100111000" => grayScale <= "00000000";
                when "100111001" => grayScale <= "00000000";
                when "100111010" => grayScale <= "00000000";
                when "100111011" => grayScale <= "00000000";
                when "101000" => grayScale <= "00000000";
                when "101001" => grayScale <= "00000000";
                when "101010" => grayScale <= "00000000";
                when "101011" => grayScale <= "00000000";
                when "1010100" => grayScale <= "00000000";
                when "1010101" => grayScale <= "00000000";
                when "1010110" => grayScale <= "00000000";
                when "1010111" => grayScale <= "00000000";
                when "10101000" => grayScale <= "00000000";
                when "10101001" => grayScale <= "00000000";
                when "10101010" => grayScale <= "00000000";
                when "10101011" => grayScale <= "00000000";
                when "10101100" => grayScale <= "00000000";
                when "10101101" => grayScale <= "00000000";
                when "10101110" => grayScale <= "00101111";
                when "10101111" => grayScale <= "01111110";
                when "101010000" => grayScale <= "01111110";
                when "101010001" => grayScale <= "01111110";
                when "101010010" => grayScale <= "00100110";
                when "101010011" => grayScale <= "00000000";
                when "101010100" => grayScale <= "00000000";
                when "101010101" => grayScale <= "00000000";
                when "101010110" => grayScale <= "00000000";
                when "101010111" => grayScale <= "00000000";
                when "101011000" => grayScale <= "00000000";
                when "101011001" => grayScale <= "00000000";
                when "101011010" => grayScale <= "00000000";
                when "101011011" => grayScale <= "00000000";
                when "101100" => grayScale <= "00000000";
                when "101101" => grayScale <= "00000000";
                when "101110" => grayScale <= "00000000";
                when "101111" => grayScale <= "00000000";
                when "1011100" => grayScale <= "00000000";
                when "1011101" => grayScale <= "00000000";
                when "1011110" => grayScale <= "00000000";
                when "1011111" => grayScale <= "00000000";
                when "10111000" => grayScale <= "00000000";
                when "10111001" => grayScale <= "00000000";
                when "10111010" => grayScale <= "00000000";
                when "10111011" => grayScale <= "00000000";
                when "10111100" => grayScale <= "00000000";
                when "10111101" => grayScale <= "00000000";
                when "10111110" => grayScale <= "01101100";
                when "10111111" => grayScale <= "01111110";
                when "101110000" => grayScale <= "01111110";
                when "101110001" => grayScale <= "01111110";
                when "101110010" => grayScale <= "00010001";
                when "101110011" => grayScale <= "00000000";
                when "101110100" => grayScale <= "00000000";
                when "101110101" => grayScale <= "00000000";
                when "101110110" => grayScale <= "00000000";
                when "101110111" => grayScale <= "00000000";
                when "101111000" => grayScale <= "00000000";
                when "101111001" => grayScale <= "00000000";
                when "101111010" => grayScale <= "00000000";
                when "101111011" => grayScale <= "00000000";
                when "110000" => grayScale <= "00000000";
                when "110001" => grayScale <= "00000000";
                when "110010" => grayScale <= "00000000";
                when "110011" => grayScale <= "00000000";
                when "1100100" => grayScale <= "00000000";
                when "1100101" => grayScale <= "00000000";
                when "1100110" => grayScale <= "00000000";
                when "1100111" => grayScale <= "00000000";
                when "11001000" => grayScale <= "00000000";
                when "11001001" => grayScale <= "00000000";
                when "11001010" => grayScale <= "00000000";
                when "11001011" => grayScale <= "00000000";
                when "11001100" => grayScale <= "00000000";
                when "11001101" => grayScale <= "00010111";
                when "11001110" => grayScale <= "01110100";
                when "11001111" => grayScale <= "01111110";
                when "110010000" => grayScale <= "01111110";
                when "110010001" => grayScale <= "00101010";
                when "110010010" => grayScale <= "00000000";
                when "110010011" => grayScale <= "00000000";
                when "110010100" => grayScale <= "00000000";
                when "110010101" => grayScale <= "00000000";
                when "110010110" => grayScale <= "00000000";
                when "110010111" => grayScale <= "00000000";
                when "110011000" => grayScale <= "00000000";
                when "110011001" => grayScale <= "00000000";
                when "110011010" => grayScale <= "00000000";
                when "110011011" => grayScale <= "00000000";
                when "110100" => grayScale <= "00000000";
                when "110101" => grayScale <= "00000000";
                when "110110" => grayScale <= "00000000";
                when "110111" => grayScale <= "00000000";
                when "1101100" => grayScale <= "00000000";
                when "1101101" => grayScale <= "00000000";
                when "1101110" => grayScale <= "00000000";
                when "1101111" => grayScale <= "00000000";
                when "11011000" => grayScale <= "00000000";
                when "11011001" => grayScale <= "00000000";
                when "11011010" => grayScale <= "00000000";
                when "11011011" => grayScale <= "00000000";
                when "11011100" => grayScale <= "00000000";
                when "11011101" => grayScale <= "01110100";
                when "11011110" => grayScale <= "01111110";
                when "11011111" => grayScale <= "01111110";
                when "110110000" => grayScale <= "01000000";
                when "110110001" => grayScale <= "00000000";
                when "110110010" => grayScale <= "00000000";
                when "110110011" => grayScale <= "00000000";
                when "110110100" => grayScale <= "00000000";
                when "110110101" => grayScale <= "00000000";
                when "110110110" => grayScale <= "00000000";
                when "110110111" => grayScale <= "00000000";
                when "110111000" => grayScale <= "00000000";
                when "110111001" => grayScale <= "00000000";
                when "110111010" => grayScale <= "00000000";
                when "110111011" => grayScale <= "00000000";
                when "111000" => grayScale <= "00000000";
                when "111001" => grayScale <= "00000000";
                when "111010" => grayScale <= "00000000";
                when "111011" => grayScale <= "00000000";
                when "1110100" => grayScale <= "00000000";
                when "1110101" => grayScale <= "00000000";
                when "1110110" => grayScale <= "00000000";
                when "1110111" => grayScale <= "00000000";
                when "11101000" => grayScale <= "00000000";
                when "11101001" => grayScale <= "00000000";
                when "11101010" => grayScale <= "00000000";
                when "11101011" => grayScale <= "00000000";
                when "11101100" => grayScale <= "00001010";
                when "11101101" => grayScale <= "01111110";
                when "11101110" => grayScale <= "01111110";
                when "11101111" => grayScale <= "01111110";
                when "111010000" => grayScale <= "00110110";
                when "111010001" => grayScale <= "00000000";
                when "111010010" => grayScale <= "00000000";
                when "111010011" => grayScale <= "00000000";
                when "111010100" => grayScale <= "00000000";
                when "111010101" => grayScale <= "00000000";
                when "111010110" => grayScale <= "00000000";
                when "111010111" => grayScale <= "00000000";
                when "111011000" => grayScale <= "00000000";
                when "111011001" => grayScale <= "00000000";
                when "111011010" => grayScale <= "00000000";
                when "111011011" => grayScale <= "00000000";
                when "111100" => grayScale <= "00000000";
                when "111101" => grayScale <= "00000000";
                when "111110" => grayScale <= "00000000";
                when "111111" => grayScale <= "00000000";
                when "1111100" => grayScale <= "00000000";
                when "1111101" => grayScale <= "00000000";
                when "1111110" => grayScale <= "00000000";
                when "1111111" => grayScale <= "00000000";
                when "11111000" => grayScale <= "00000000";
                when "11111001" => grayScale <= "00000000";
                when "11111010" => grayScale <= "00000000";
                when "11111011" => grayScale <= "00001010";
                when "11111100" => grayScale <= "01100111";
                when "11111101" => grayScale <= "01111110";
                when "11111110" => grayScale <= "01111110";
                when "11111111" => grayScale <= "01110011";
                when "111110000" => grayScale <= "00010111";
                when "111110001" => grayScale <= "00000000";
                when "111110010" => grayScale <= "00000000";
                when "111110011" => grayScale <= "00000000";
                when "111110100" => grayScale <= "00000000";
                when "111110101" => grayScale <= "00000000";
                when "111110110" => grayScale <= "00000000";
                when "111110111" => grayScale <= "00000000";
                when "111111000" => grayScale <= "00000000";
                when "111111001" => grayScale <= "00000000";
                when "111111010" => grayScale <= "00000000";
                when "111111011" => grayScale <= "00000000";
                when "1000000" => grayScale <= "00000000";
                when "1000001" => grayScale <= "00000000";
                when "1000010" => grayScale <= "00000000";
                when "1000011" => grayScale <= "00000000";
                when "10000100" => grayScale <= "00000000";
                when "10000101" => grayScale <= "00000000";
                when "10000110" => grayScale <= "00000000";
                when "10000111" => grayScale <= "00000000";
                when "100001000" => grayScale <= "00000000";
                when "100001001" => grayScale <= "00000000";
                when "100001010" => grayScale <= "00000000";
                when "100001011" => grayScale <= "01011011";
                when "100001100" => grayScale <= "01111110";
                when "100001101" => grayScale <= "10000000";
                when "100001110" => grayScale <= "01101111";
                when "100001111" => grayScale <= "00010100";
                when "1000010000" => grayScale <= "00000000";
                when "1000010001" => grayScale <= "00000000";
                when "1000010010" => grayScale <= "00000000";
                when "1000010011" => grayScale <= "00000000";
                when "1000010100" => grayScale <= "00000000";
                when "1000010101" => grayScale <= "00000000";
                when "1000010110" => grayScale <= "00000000";
                when "1000010111" => grayScale <= "00000000";
                when "1000011000" => grayScale <= "00000000";
                when "1000011001" => grayScale <= "00000000";
                when "1000011010" => grayScale <= "00000000";
                when "1000011011" => grayScale <= "00000000";
                when "1000100" => grayScale <= "00000000";
                when "1000101" => grayScale <= "00000000";
                when "1000110" => grayScale <= "00000000";
                when "1000111" => grayScale <= "00000000";
                when "10001100" => grayScale <= "00000000";
                when "10001101" => grayScale <= "00000000";
                when "10001110" => grayScale <= "00000000";
                when "10001111" => grayScale <= "00000000";
                when "100011000" => grayScale <= "00000000";
                when "100011001" => grayScale <= "00000000";
                when "100011010" => grayScale <= "00001010";
                when "100011011" => grayScale <= "01100100";
                when "100011100" => grayScale <= "01111110";
                when "100011101" => grayScale <= "01111110";
                when "100011110" => grayScale <= "01011001";
                when "100011111" => grayScale <= "00000000";
                when "1000110000" => grayScale <= "00000000";
                when "1000110001" => grayScale <= "00000000";
                when "1000110010" => grayScale <= "00000000";
                when "1000110011" => grayScale <= "00000000";
                when "1000110100" => grayScale <= "00000000";
                when "1000110101" => grayScale <= "00000000";
                when "1000110110" => grayScale <= "00000000";
                when "1000110111" => grayScale <= "00000000";
                when "1000111000" => grayScale <= "00000000";
                when "1000111001" => grayScale <= "00000000";
                when "1000111010" => grayScale <= "00000000";
                when "1000111011" => grayScale <= "00000000";
                when "1001000" => grayScale <= "00000000";
                when "1001001" => grayScale <= "00000000";
                when "1001010" => grayScale <= "00000000";
                when "1001011" => grayScale <= "00000000";
                when "10010100" => grayScale <= "00000000";
                when "10010101" => grayScale <= "00000000";
                when "10010110" => grayScale <= "00000000";
                when "10010111" => grayScale <= "00000000";
                when "100101000" => grayScale <= "00000000";
                when "100101001" => grayScale <= "00001000";
                when "100101010" => grayScale <= "00110001";
                when "100101011" => grayScale <= "01111110";
                when "100101100" => grayScale <= "01111110";
                when "100101101" => grayScale <= "01111110";
                when "100101110" => grayScale <= "00100110";
                when "100101111" => grayScale <= "00000000";
                when "1001010000" => grayScale <= "00000000";
                when "1001010001" => grayScale <= "00000000";
                when "1001010010" => grayScale <= "00000000";
                when "1001010011" => grayScale <= "00000000";
                when "1001010100" => grayScale <= "00000000";
                when "1001010101" => grayScale <= "00000000";
                when "1001010110" => grayScale <= "00000000";
                when "1001010111" => grayScale <= "00000000";
                when "1001011000" => grayScale <= "00000000";
                when "1001011001" => grayScale <= "00000000";
                when "1001011010" => grayScale <= "00000000";
                when "1001011011" => grayScale <= "00000000";
                when "1001100" => grayScale <= "00000000";
                when "1001101" => grayScale <= "00000000";
                when "1001110" => grayScale <= "00000000";
                when "1001111" => grayScale <= "00000000";
                when "10011100" => grayScale <= "00000000";
                when "10011101" => grayScale <= "00000000";
                when "10011110" => grayScale <= "00000000";
                when "10011111" => grayScale <= "00000000";
                when "100111000" => grayScale <= "00000000";
                when "100111001" => grayScale <= "00110110";
                when "100111010" => grayScale <= "01111110";
                when "100111011" => grayScale <= "01111110";
                when "100111100" => grayScale <= "01111110";
                when "100111101" => grayScale <= "01011111";
                when "100111110" => grayScale <= "00000111";
                when "100111111" => grayScale <= "00000000";
                when "1001110000" => grayScale <= "00000000";
                when "1001110001" => grayScale <= "00000000";
                when "1001110010" => grayScale <= "00000000";
                when "1001110011" => grayScale <= "00000000";
                when "1001110100" => grayScale <= "00000000";
                when "1001110101" => grayScale <= "00000000";
                when "1001110110" => grayScale <= "00000000";
                when "1001110111" => grayScale <= "00000000";
                when "1001111000" => grayScale <= "00000000";
                when "1001111001" => grayScale <= "00000000";
                when "1001111010" => grayScale <= "00000000";
                when "1001111011" => grayScale <= "00000000";
                when "1010000" => grayScale <= "00000000";
                when "1010001" => grayScale <= "00000000";
                when "1010010" => grayScale <= "00000000";
                when "1010011" => grayScale <= "00000000";
                when "10100100" => grayScale <= "00000000";
                when "10100101" => grayScale <= "00000000";
                when "10100110" => grayScale <= "00000000";
                when "10100111" => grayScale <= "00000000";
                when "101001000" => grayScale <= "00000000";
                when "101001001" => grayScale <= "01010101";
                when "101001010" => grayScale <= "01111110";
                when "101001011" => grayScale <= "01111110";
                when "101001100" => grayScale <= "01111110";
                when "101001101" => grayScale <= "00000000";
                when "101001110" => grayScale <= "00000000";
                when "101001111" => grayScale <= "00000000";
                when "1010010000" => grayScale <= "00000000";
                when "1010010001" => grayScale <= "00000000";
                when "1010010010" => grayScale <= "00000000";
                when "1010010011" => grayScale <= "00000000";
                when "1010010100" => grayScale <= "00000000";
                when "1010010101" => grayScale <= "00000000";
                when "1010010110" => grayScale <= "00000000";
                when "1010010111" => grayScale <= "00000000";
                when "1010011000" => grayScale <= "00000000";
                when "1010011001" => grayScale <= "00000000";
                when "1010011010" => grayScale <= "00000000";
                when "1010011011" => grayScale <= "00000000";
                when "1010100" => grayScale <= "00000000";
                when "1010101" => grayScale <= "00000000";
                when "1010110" => grayScale <= "00000000";
                when "1010111" => grayScale <= "00000000";
                when "10101100" => grayScale <= "00000000";
                when "10101101" => grayScale <= "00000000";
                when "10101110" => grayScale <= "00000000";
                when "10101111" => grayScale <= "00000000";
                when "101011000" => grayScale <= "00010101";
                when "101011001" => grayScale <= "01111110";
                when "101011010" => grayScale <= "01111110";
                when "101011011" => grayScale <= "01111110";
                when "101011100" => grayScale <= "01111110";
                when "101011101" => grayScale <= "00000000";
                when "101011110" => grayScale <= "00000000";
                when "101011111" => grayScale <= "00000000";
                when "1010110000" => grayScale <= "00000000";
                when "1010110001" => grayScale <= "00000000";
                when "1010110010" => grayScale <= "00000000";
                when "1010110011" => grayScale <= "00000000";
                when "1010110100" => grayScale <= "00000000";
                when "1010110101" => grayScale <= "00000000";
                when "1010110110" => grayScale <= "00000000";
                when "1010110111" => grayScale <= "00000000";
                when "1010111000" => grayScale <= "00000000";
                when "1010111001" => grayScale <= "00000000";
                when "1010111010" => grayScale <= "00000000";
                when "1010111011" => grayScale <= "00000000";
                when "1011000" => grayScale <= "00000000";
                when "1011001" => grayScale <= "00000000";
                when "1011010" => grayScale <= "00000000";
                when "1011011" => grayScale <= "00000000";
                when "10110100" => grayScale <= "00000000";
                when "10110101" => grayScale <= "00000000";
                when "10110110" => grayScale <= "00000000";
                when "10110111" => grayScale <= "00000000";
                when "101101000" => grayScale <= "00111110";
                when "101101001" => grayScale <= "01111110";
                when "101101010" => grayScale <= "01111110";
                when "101101011" => grayScale <= "01111110";
                when "101101100" => grayScale <= "01111110";
                when "101101101" => grayScale <= "00110100";
                when "101101110" => grayScale <= "00000000";
                when "101101111" => grayScale <= "00000000";
                when "1011010000" => grayScale <= "00000000";
                when "1011010001" => grayScale <= "00000000";
                when "1011010010" => grayScale <= "00000000";
                when "1011010011" => grayScale <= "00000000";
                when "1011010100" => grayScale <= "00000000";
                when "1011010101" => grayScale <= "00000000";
                when "1011010110" => grayScale <= "00000000";
                when "1011010111" => grayScale <= "00000000";
                when "1011011000" => grayScale <= "00000000";
                when "1011011001" => grayScale <= "00000000";
                when "1011011010" => grayScale <= "00000000";
                when "1011011011" => grayScale <= "00000000";
                when "1011100" => grayScale <= "00000000";
                when "1011101" => grayScale <= "00000000";
                when "1011110" => grayScale <= "00000000";
                when "1011111" => grayScale <= "00000000";
                when "10111100" => grayScale <= "00000000";
                when "10111101" => grayScale <= "00000000";
                when "10111110" => grayScale <= "00000000";
                when "10111111" => grayScale <= "00000000";
                when "101111000" => grayScale <= "00000000";
                when "101111001" => grayScale <= "01010100";
                when "101111010" => grayScale <= "01111110";
                when "101111011" => grayScale <= "01111110";
                when "101111100" => grayScale <= "01111110";
                when "101111101" => grayScale <= "00011111";
                when "101111110" => grayScale <= "00000000";
                when "101111111" => grayScale <= "00000000";
                when "1011110000" => grayScale <= "00000000";
                when "1011110001" => grayScale <= "00000000";
                when "1011110010" => grayScale <= "00000000";
                when "1011110011" => grayScale <= "00000000";
                when "1011110100" => grayScale <= "00000000";
                when "1011110101" => grayScale <= "00000000";
                when "1011110110" => grayScale <= "00000000";
                when "1011110111" => grayScale <= "00000000";
                when "1011111000" => grayScale <= "00000000";
                when "1011111001" => grayScale <= "00000000";
                when "1011111010" => grayScale <= "00000000";
                when "1011111011" => grayScale <= "00000000";
                when "1100000" => grayScale <= "00000000";
                when "1100001" => grayScale <= "00000000";
                when "1100010" => grayScale <= "00000000";
                when "1100011" => grayScale <= "00000000";
                when "11000100" => grayScale <= "00000000";
                when "11000101" => grayScale <= "00000000";
                when "11000110" => grayScale <= "00000000";
                when "11000111" => grayScale <= "00000000";
                when "110001000" => grayScale <= "00000000";
                when "110001001" => grayScale <= "00000000";
                when "110001010" => grayScale <= "00000000";
                when "110001011" => grayScale <= "00000000";
                when "110001100" => grayScale <= "00000000";
                when "110001101" => grayScale <= "00000000";
                when "110001110" => grayScale <= "00000000";
                when "110001111" => grayScale <= "00000000";
                when "1100010000" => grayScale <= "00000000";
                when "1100010001" => grayScale <= "00000000";
                when "1100010010" => grayScale <= "00000000";
                when "1100010011" => grayScale <= "00000000";
                when "1100010100" => grayScale <= "00000000";
                when "1100010101" => grayScale <= "00000000";
                when "1100010110" => grayScale <= "00000000";
                when "1100010111" => grayScale <= "00000000";
                when "1100011000" => grayScale <= "00000000";
                when "1100011001" => grayScale <= "00000000";
                when "1100011010" => grayScale <= "00000000";
                when "1100011011" => grayScale <= "00000000";
                when "1100100" => grayScale <= "00000000";
                when "1100101" => grayScale <= "00000000";
                when "1100110" => grayScale <= "00000000";
                when "1100111" => grayScale <= "00000000";
                when "11001100" => grayScale <= "00000000";
                when "11001101" => grayScale <= "00000000";
                when "11001110" => grayScale <= "00000000";
                when "11001111" => grayScale <= "00000000";
                when "110011000" => grayScale <= "00000000";
                when "110011001" => grayScale <= "00000000";
                when "110011010" => grayScale <= "00000000";
                when "110011011" => grayScale <= "00000000";
                when "110011100" => grayScale <= "00000000";
                when "110011101" => grayScale <= "00000000";
                when "110011110" => grayScale <= "00000000";
                when "110011111" => grayScale <= "00000000";
                when "1100110000" => grayScale <= "00000000";
                when "1100110001" => grayScale <= "00000000";
                when "1100110010" => grayScale <= "00000000";
                when "1100110011" => grayScale <= "00000000";
                when "1100110100" => grayScale <= "00000000";
                when "1100110101" => grayScale <= "00000000";
                when "1100110110" => grayScale <= "00000000";
                when "1100110111" => grayScale <= "00000000";
                when "1100111000" => grayScale <= "00000000";
                when "1100111001" => grayScale <= "00000000";
                when "1100111010" => grayScale <= "00000000";
                when "1100111011" => grayScale <= "00000000";
                when "1101000" => grayScale <= "00000000";
                when "1101001" => grayScale <= "00000000";
                when "1101010" => grayScale <= "00000000";
                when "1101011" => grayScale <= "00000000";
                when "11010100" => grayScale <= "00000000";
                when "11010101" => grayScale <= "00000000";
                when "11010110" => grayScale <= "00000000";
                when "11010111" => grayScale <= "00000000";
                when "110101000" => grayScale <= "00000000";
                when "110101001" => grayScale <= "00000000";
                when "110101010" => grayScale <= "00000000";
                when "110101011" => grayScale <= "00000000";
                when "110101100" => grayScale <= "00000000";
                when "110101101" => grayScale <= "00000000";
                when "110101110" => grayScale <= "00000000";
                when "110101111" => grayScale <= "00000000";
                when "1101010000" => grayScale <= "00000000";
                when "1101010001" => grayScale <= "00000000";
                when "1101010010" => grayScale <= "00000000";
                when "1101010011" => grayScale <= "00000000";
                when "1101010100" => grayScale <= "00000000";
                when "1101010101" => grayScale <= "00000000";
                when "1101010110" => grayScale <= "00000000";
                when "1101010111" => grayScale <= "00000000";
                when "1101011000" => grayScale <= "00000000";
                when "1101011001" => grayScale <= "00000000";
                when "1101011010" => grayScale <= "00000000";
                when "1101011011" => grayScale <= "00000000";
                when "1101100" => grayScale <= "00000000";
                when "1101101" => grayScale <= "00000000";
                when "1101110" => grayScale <= "00000000";
                when "1101111" => grayScale <= "00000000";
                when "11011100" => grayScale <= "00000000";
                when "11011101" => grayScale <= "00000000";
                when "11011110" => grayScale <= "00000000";
                when "11011111" => grayScale <= "00000000";
                when "110111000" => grayScale <= "00000000";
                when "110111001" => grayScale <= "00000000";
                when "110111010" => grayScale <= "00000000";
                when "110111011" => grayScale <= "00000000";
                when "110111100" => grayScale <= "00000000";
                when "110111101" => grayScale <= "00000000";
                when "110111110" => grayScale <= "00000000";
                when "110111111" => grayScale <= "00000000";
                when "1101110000" => grayScale <= "00000000";
                when "1101110001" => grayScale <= "00000000";
                when "1101110010" => grayScale <= "00000000";
                when "1101110011" => grayScale <= "00000000";
                when "1101110100" => grayScale <= "00000000";
                when "1101110101" => grayScale <= "00000000";
                when "1101110110" => grayScale <= "00000000";
                when "1101110111" => grayScale <= "00000000";
                when "1101111000" => grayScale <= "00000000";
                when "1101111001" => grayScale <= "00000000";
                when "1101111010" => grayScale <= "00000000";
                when "1101111011" => grayScale <= "00000000";
                when others => grayScale <= "00000000";
        end case;
    end if;
    end process;
end;
